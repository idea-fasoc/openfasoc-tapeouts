** sch_path:
*+ /home/andylithia/openmpw/openfasoc-tapeouts/gf180mcu_padframe/tb/digital_io_switching.sch
**.subckt digital_io_switching
V1 DVDD GND 3
.save i(v1)
V2 VDD GND 3
.save i(v2)
V3 DVSS GND 0
.save i(v3)
V4 VSS GND 0
.save i(v4)
V5 A GND PULSE(0 3 10n 100p 100p 10n 20n)
.save i(v5)
V6 PDRV1 GND 3
.save i(v6)
V7 IE GND 3
.save i(v7)
V8 OE GND 3
.save i(v8)
V9 PU GND 0
.save i(v9)
V10 PD GND 0
.save i(v10)
V11 SL GND 0
.save i(v11)
V12 PDRV0 GND 3
.save i(v12)
V13 CS GND 3.3
.save i(v13)
**** begin user architecture code


.tran 100p 100n
.save all
.control
run
display
plot A PAD0 Y0
plot PAD0 PAD1 PAD2 PAD3
.endc



.include /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice diode_typical
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical


.include ../gf180mcu_fd_io.spice
XDUT0 A CS DVDD DVSS IE OE PAD0 PD VSS VSS PU SL VDD VSS Y0 gf180mcu_fd_io__bi_t
XDUT1 A CS DVDD DVSS IE OE PAD1 PD VDD VSS PU SL VDD VSS Y1 gf180mcu_fd_io__bi_t
XDUT2 A CS DVDD DVSS IE OE PAD2 PD VSS VDD PU SL VDD VSS Y2 gf180mcu_fd_io__bi_t
XDUT3 A CS DVDD DVSS IE OE PAD3 PD VDD VDD PU SL VDD VSS Y3 gf180mcu_fd_io__bi_t

**** end user architecture code
**.ends
.GLOBAL GND
.end
