** sch_path: /home/andylithia/openmpw/openfasoc-tapeouts/gf180mcu_padframe/tb/analog_io_sppex.sch
**.subckt analog_io_sppex
V1 DVDD GND 3
.save i(v1)
V2 VDD GND 3
.save i(v2)
V3 DVSS GND 0
.save i(v3)
V4 VSS GND 0
.save i(v4)
V5 net1 GND DC 3 AC 1
.save i(v5)
R1 ASIG net1 1k m=1
**** begin user architecture code


.ac dec 100 1k 100G
.save all
.control
run
display
plot PAD ASIG
plot vdb(asig) vdb(pad)
.endc



.include /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice diode_typical
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical
.lib /home/andylithia/openmpw/pdk_1/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical


.include ./gf180mcu_fd_io__asig_5p0_extracted.spice
XDUT DVSS DVDD VSS VDD PAD ASIG gf180mcu_fd_io__asig_5p0_extracted

**** end user architecture code
**.ends
.GLOBAL GND
.end
