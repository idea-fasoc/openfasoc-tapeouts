.subckt gf180mcu_fd_io__asig_5p0_extracted  DVSS DVDD VSS VDD PAD ASIG5V
cDVDD/0 DVDD:16209 vss 7.57208f
cDVDD/1 DVDD:16205 vss 79.679f
cDVDD/2 DVDD:16160 vss 7.5076f
cDVDD/3 DVDD:16156 vss 78.2189f
cDVDD/4 DVDD:16083 vss 20.7374f
cDVDD/5 DVDD:15976 vss 21.0976f
cDVDD/6 DVDD:15870 vss 20.8618f
cDVDD/7 DVDD:15757 vss 0.56211f
cDVDD/8 DVDD:15753 vss 0.581688f
cDVDD/9 DVDD:15743 vss 0.221594f
cDVDD/10 DVDD:15733 vss 0.1849f
cDVDD/11 DVDD:15724 vss 0.526184f
cDVDD/12 DVDD:15714 vss 0.26583f
cDVDD/13 DVDD:15704 vss 0.303359f
cDVDD/14 DVDD:15695 vss 2.74937f
cDVDD/15 DVDD:15691 vss 0.101053f
cDVDD/16 DVDD:15686 vss 0.457353f
cDVDD/17 DVDD:15677 vss 14.1501f
cDVDD/18 DVDD:15468 vss 28.2397f
cDVDD/19 DVDD:15436 vss 202.45f
cDVDD/20 DVDD:15435 vss 5.38399f
cDVDD/21 DVDD:15426 vss 33.6478f
cDVDD/22 DVDD:15416 vss 16.376f
cDVDD/23 DVDD:15412 vss 1.61205f
cDVDD/24 DVDD:15373 vss 23.1914f
cDVDD/25 DVDD:15295 vss 17.1363f
cDVDD/26 DVDD:15004 vss 32.7136f
cDVDD/27 DVDD:14722 vss 26.6155f
cDVDD/28 DVDD:14437 vss 26.6155f
cDVDD/29 DVDD:14155 vss 32.7132f
cDVDD/30 DVDD:14082 vss 16.468f
cDVDD/31 DVDD:14078 vss 1.62203f
cDVDD/32 DVDD:14039 vss 23.4037f
cDVDD/33 DVDD:13961 vss 17.1363f
cDVDD/34 DVDD:13695 vss 1.19876f
cDVDD/35 DVDD:13645 vss 2.93002f
cDVDD/36 DVDD:13626 vss 3.93797f
cDVDD/37 DVDD:13607 vss 3.46682f
cDVDD/38 DVDD:13599 vss 1.17601f
cDVDD/39 DVDD:13432 vss 31.9204f
cDVDD/40 DVDD:13120 vss 36.606f
cDVDD/41 DVDD:12805 vss 30.0321f
cDVDD/42 DVDD:12490 vss 30.0321f
cDVDD/43 DVDD:12069 vss 36.6052f
cDVDD/44 DVDD:11910 vss 6.35693f
cDVDD/45 DVDD:11814 vss 6.45956f
cDVDD/46 DVDD:11718 vss 6.45956f
cDVDD/47 DVDD:11622 vss 6.35822f
cDVDD/48 DVDD:11300 vss 16.3982f
cDVDD/49 DVDD:11280 vss 0.60798f
cDVDD/50 DVDD:11228 vss 2.20998f
cDVDD/51 DVDD:11223 vss 0.246528f
cDVDD/52 DVDD:11183 vss 2.61894f
cDVDD/53 DVDD:11175 vss 0.283361f
cDVDD/54 DVDD:11149 vss 12.246f
cDVDD/55 DVDD:11112 vss 12.276f
cDVDD/56 DVDD:11080 vss 8.21533f
cDVDD/57 DVDD vss 13.7761f
cDVDD/58 DVDD:11060 vss 16.7658f
cDVDD/59 DVDD:11056 vss 10.008f
cDVDD/60 DVDD:10963 vss 16.9075f
cDVDD/61 DVDD:10959 vss 10.0118f
cDVDD/62 DVDD:10866 vss 16.7995f
cDVDD/63 DVDD:10862 vss 10.002f
cDVDD/64 DVDD:10771 vss 0.18771f
cDVDD/65 DVDD:10766 vss 0.314239f
cDVDD/66 DVDD:10761 vss 0.675686f
cDVDD/67 DVDD:10757 vss 0.20557f
cDVDD/68 DVDD:10752 vss 0.205558f
cDVDD/69 DVDD:10727 vss 1.00758f
cDVDD/70 DVDD:10717 vss 1.00236f
cDVDD/71 DVDD:10688 vss 3.72855f
cDVDD/72 DVDD:10683 vss 0.197672f
cDVDD/73 DVDD:10663 vss 2.33273f
cDVDD/74 DVDD:10658 vss 0.193915f
cDVDD/75 D8:neg vss 0.845741f
cDVDD/76 DVDD:9148 vss 0.459122f
cDVDD/77 DVDD:9140 vss 12.6303f
cDVDD/78 DVDD:9133 vss 2.45177f
cDVDD/79 DVDD:9125 vss 2.42021f
cDVDD/80 DVDD:9116 vss 0.607574f
cDVDD/81 X52/X1/X2/X1/C0:pos vss 4.1609f
cDVDD/82 DVDD:9086 vss 0.058323f
cDVDD/83 DVDD:9078 vss 16.9289f
cDVDD/84 DVDD:9071 vss 2.39888f
cDVDD/85 DVDD:9063 vss 2.44184f
cDVDD/86 DVDD:9054 vss 0.0771812f
cDVDD/87 X52/X1/X2/X0/C0:pos vss 4.95726f
cDVDD/88 DVDD:8976 vss 0.058323f
cDVDD/89 DVDD:8968 vss 16.9289f
cDVDD/90 DVDD:8961 vss 2.39888f
cDVDD/91 DVDD:8953 vss 2.44184f
cDVDD/92 DVDD:8944 vss 0.0771812f
cDVDD/93 X52/X1/X1/X1/C0:pos vss 4.95726f
cDVDD/94 DVDD:8906 vss 14.3793f
cDVDD/95 DVDD:8899 vss 2.39421f
cDVDD/96 DVDD:8891 vss 2.42622f
cDVDD/97 X52/X1/X1/X0/C0:pos vss 4.20338f
cDVDD/98 DVDD:8698 vss 0.457738f
cDVDD/99 DVDD:8690 vss 12.4577f
cDVDD/100 DVDD:8683 vss 2.39209f
cDVDD/101 DVDD:8675 vss 2.42019f
cDVDD/102 DVDD:8666 vss 0.605744f
cDVDD/103 X52/X0/X2/X1/C0:pos vss 4.16126f
cDVDD/104 DVDD:8636 vss 0.0568369f
cDVDD/105 DVDD:8628 vss 16.7695f
cDVDD/106 DVDD:8621 vss 2.3988f
cDVDD/107 DVDD:8613 vss 2.44179f
cDVDD/108 DVDD:8604 vss 0.0752146f
cDVDD/109 X52/X0/X2/X0/C0:pos vss 4.95799f
cDVDD/110 DVDD:8526 vss 0.0568369f
cDVDD/111 DVDD:8518 vss 16.7695f
cDVDD/112 DVDD:8511 vss 2.3988f
cDVDD/113 DVDD:8503 vss 2.44179f
cDVDD/114 DVDD:8494 vss 0.0752146f
cDVDD/115 X52/X0/X1/X1/C0:pos vss 4.95799f
cDVDD/116 DVDD:8456 vss 14.4709f
cDVDD/117 DVDD:8449 vss 2.39809f
cDVDD/118 DVDD:8441 vss 2.42619f
cDVDD/119 X52/X0/X1/X0/C0:pos vss 4.20791f
cDVDD/120 DVDD:8104 vss 0.457289f
cDVDD/121 DVDD:8096 vss 12.2929f
cDVDD/122 DVDD:8089 vss 2.39213f
cDVDD/123 DVDD:8081 vss 2.40438f
cDVDD/124 DVDD:8072 vss 0.605149f
cDVDD/125 X51/X1/X2/X1/C0:pos vss 4.16073f
cDVDD/126 DVDD:8042 vss 0.056491f
cDVDD/127 DVDD:8034 vss 16.636f
cDVDD/128 DVDD:8027 vss 2.39888f
cDVDD/129 DVDD:8019 vss 2.43633f
cDVDD/130 DVDD:8010 vss 0.0747568f
cDVDD/131 X51/X1/X2/X0/C0:pos vss 4.95687f
cDVDD/132 DVDD:7932 vss 0.056491f
cDVDD/133 DVDD:7924 vss 16.636f
cDVDD/134 DVDD:7917 vss 2.39888f
cDVDD/135 DVDD:7909 vss 2.43633f
cDVDD/136 DVDD:7900 vss 0.0747568f
cDVDD/137 X51/X1/X1/X1/C0:pos vss 4.95687f
cDVDD/138 DVDD:7862 vss 14.3236f
cDVDD/139 DVDD:7855 vss 2.39813f
cDVDD/140 DVDD:7847 vss 2.41038f
cDVDD/141 X51/X1/X1/X0/C0:pos vss 4.20739f
cDVDD/142 DVDD:7654 vss 0.455658f
cDVDD/143 DVDD:7646 vss 12.541f
cDVDD/144 DVDD:7639 vss 2.39209f
cDVDD/145 DVDD:7631 vss 2.40438f
cDVDD/146 DVDD:7622 vss 0.602991f
cDVDD/147 X51/X0/X2/X1/C0:pos vss 4.16126f
cDVDD/148 DVDD:7592 vss 0.0547567f
cDVDD/149 DVDD:7584 vss 16.8412f
cDVDD/150 DVDD:7577 vss 2.3988f
cDVDD/151 DVDD:7569 vss 2.43633f
cDVDD/152 DVDD:7560 vss 0.0724618f
cDVDD/153 X51/X0/X2/X0/C0:pos vss 4.95798f
cDVDD/154 DVDD:7482 vss 0.0547567f
cDVDD/155 DVDD:7474 vss 16.8412f
cDVDD/156 DVDD:7467 vss 2.3988f
cDVDD/157 DVDD:7459 vss 2.43633f
cDVDD/158 DVDD:7450 vss 0.0724618f
cDVDD/159 X51/X0/X1/X1/C0:pos vss 4.95798f
cDVDD/160 DVDD:7412 vss 14.4612f
cDVDD/161 DVDD:7405 vss 2.39809f
cDVDD/162 DVDD:7397 vss 2.40362f
cDVDD/163 X51/X0/X1/X0/C0:pos vss 4.20829f
cDVDD/164 DVDD:7060 vss 0.459993f
cDVDD/165 DVDD:7052 vss 12.663f
cDVDD/166 DVDD:7045 vss 2.39209f
cDVDD/167 DVDD:7037 vss 2.40979f
cDVDD/168 DVDD:7028 vss 0.608728f
cDVDD/169 X50/X1/X2/X1/C0:pos vss 4.1609f
cDVDD/170 DVDD:6998 vss 0.0590918f
cDVDD/171 DVDD:6990 vss 16.9175f
cDVDD/172 DVDD:6983 vss 2.3988f
cDVDD/173 DVDD:6975 vss 2.43633f
cDVDD/174 DVDD:6966 vss 0.0781985f
cDVDD/175 X50/X1/X2/X0/C0:pos vss 4.95727f
cDVDD/176 DVDD:6888 vss 0.0590918f
cDVDD/177 DVDD:6880 vss 16.9175f
cDVDD/178 DVDD:6873 vss 2.3988f
cDVDD/179 DVDD:6865 vss 2.44121f
cDVDD/180 DVDD:6856 vss 0.0781985f
cDVDD/181 X50/X1/X1/X1/C0:pos vss 4.95727f
cDVDD/182 DVDD:6818 vss 13.9735f
cDVDD/183 DVDD:6811 vss 2.39422f
cDVDD/184 DVDD:6803 vss 2.40359f
cDVDD/185 X50/X1/X1/X0/C0:pos vss 4.19337f
cDVDD/186 DVDD:6610 vss 0.455658f
cDVDD/187 DVDD:6602 vss 12.296f
cDVDD/188 DVDD:6595 vss 2.39752f
cDVDD/189 DVDD:6587 vss 2.40979f
cDVDD/190 DVDD:6578 vss 0.602991f
cDVDD/191 X50/X0/X2/X1/C0:pos vss 4.16054f
cDVDD/192 DVDD:6548 vss 0.0547567f
cDVDD/193 DVDD:6540 vss 16.6032f
cDVDD/194 DVDD:6533 vss 2.40613f
cDVDD/195 DVDD:6525 vss 2.43633f
cDVDD/196 DVDD:6516 vss 0.0724618f
cDVDD/197 X50/X0/X2/X0/C0:pos vss 4.95654f
cDVDD/198 DVDD:6438 vss 0.0547567f
cDVDD/199 DVDD:6430 vss 16.6032f
cDVDD/200 DVDD:6423 vss 2.40429f
cDVDD/201 DVDD:6415 vss 2.44121f
cDVDD/202 DVDD:6406 vss 0.0724618f
cDVDD/203 X50/X0/X1/X1/C0:pos vss 4.95654f
cDVDD/204 DVDD:6368 vss 13.4264f
cDVDD/205 DVDD:6361 vss 2.40119f
cDVDD/206 DVDD:6353 vss 2.40979f
cDVDD/207 X50/X0/X1/X0/C0:pos vss 4.16355f
cDVDD/208 DVDD:6016 vss 0.458129f
cDVDD/209 DVDD:6008 vss 12.5082f
cDVDD/210 DVDD:6001 vss 2.40119f
cDVDD/211 DVDD:5993 vss 2.40979f
cDVDD/212 DVDD:5984 vss 0.606261f
cDVDD/213 X49/X1/X2/X1/C0:pos vss 4.16126f
cDVDD/214 DVDD:5954 vss 0.0572278f
cDVDD/215 DVDD:5946 vss 16.7737f
cDVDD/216 DVDD:5939 vss 2.40613f
cDVDD/217 DVDD:5931 vss 2.43633f
cDVDD/218 DVDD:5922 vss 0.0757318f
cDVDD/219 X49/X1/X2/X0/C0:pos vss 4.95794f
cDVDD/220 DVDD:5844 vss 0.0572278f
cDVDD/221 DVDD:5836 vss 16.7737f
cDVDD/222 DVDD:5829 vss 2.40429f
cDVDD/223 DVDD:5821 vss 2.44121f
cDVDD/224 DVDD:5812 vss 0.0757318f
cDVDD/225 X49/X1/X1/X1/C0:pos vss 4.95794f
cDVDD/226 DVDD:5774 vss 13.7264f
cDVDD/227 DVDD:5767 vss 2.40119f
cDVDD/228 DVDD:5759 vss 2.40979f
cDVDD/229 X49/X1/X1/X0/C0:pos vss 4.18159f
cDVDD/230 DVDD:5566 vss 0.455658f
cDVDD/231 DVDD:5558 vss 12.2936f
cDVDD/232 DVDD:5551 vss 2.40119f
cDVDD/233 DVDD:5543 vss 2.40762f
cDVDD/234 DVDD:5534 vss 0.602991f
cDVDD/235 X49/X0/X2/X1/C0:pos vss 4.16054f
cDVDD/236 DVDD:5504 vss 0.0547567f
cDVDD/237 DVDD:5496 vss 16.5989f
cDVDD/238 DVDD:5489 vss 2.40796f
cDVDD/239 DVDD:5481 vss 2.43417f
cDVDD/240 DVDD:5472 vss 0.0724618f
cDVDD/241 X49/X0/X2/X0/C0:pos vss 4.95654f
cDVDD/242 DVDD:5394 vss 0.0547567f
cDVDD/243 DVDD:5386 vss 16.5989f
cDVDD/244 DVDD:5379 vss 2.40613f
cDVDD/245 DVDD:5371 vss 2.44391f
cDVDD/246 DVDD:5362 vss 0.0724618f
cDVDD/247 X49/X0/X1/X1/C0:pos vss 4.95654f
cDVDD/248 DVDD:5324 vss 13.4269f
cDVDD/249 DVDD:5317 vss 2.40119f
cDVDD/250 DVDD:5309 vss 2.40762f
cDVDD/251 X49/X0/X1/X0/C0:pos vss 4.16349f
cDVDD/252 DVDD:5116 vss 0.391353f
cDVDD/253 DVDD:5108 vss 12.6482f
cDVDD/254 DVDD:5101 vss 2.38986f
cDVDD/255 DVDD:5093 vss 2.42012f
cDVDD/256 DVDD:5084 vss 0.517893f
cDVDD/257 X48/X2/X1/C0:pos vss 4.16124f
cDVDD/258 DVDD:5054 vss 0.0568369f
cDVDD/259 DVDD:5046 vss 16.7651f
cDVDD/260 DVDD:5039 vss 2.39663f
cDVDD/261 DVDD:5031 vss 2.44179f
cDVDD/262 DVDD:5022 vss 0.0752146f
cDVDD/263 X48/X2/X0/C0:pos vss 4.95799f
cDVDD/264 DVDD:4944 vss 0.0568369f
cDVDD/265 DVDD:4936 vss 16.7651f
cDVDD/266 DVDD:4929 vss 2.39663f
cDVDD/267 DVDD:4921 vss 2.44179f
cDVDD/268 DVDD:4912 vss 0.0752146f
cDVDD/269 X48/X1/X1/C0:pos vss 4.95799f
cDVDD/270 DVDD:4874 vss 13.8491f
cDVDD/271 DVDD:4867 vss 2.39465f
cDVDD/272 DVDD:4859 vss 2.42548f
cDVDD/273 X48/X1/X0/C0:pos vss 4.17947f
cDVDD/274 DVDD:4222 vss 0.413659f
cDVDD/275 DVDD:4221 vss 33.0042f
cDVDD/276 DVDD:4212 vss 0.363814f
cDVDD/277 DVDD:4202 vss 0.363814f
cDVDD/278 DVDD:4192 vss 0.363814f
cDVDD/279 DVDD:4182 vss 4.26589f
cDVDD/280 DVDD:4178 vss 7.88579f
cDVDD/281 DVDD:4174 vss 7.89665f
cDVDD/282 DVDD:4170 vss 7.88579f
cDVDD/283 DVDD:4168 vss 3.14615f
cDVDD/284 DVDD:4165 vss 37.1713f
cDVDD/285 DVDD:4133 vss 37.308f
cDVDD/286 DVDD:4101 vss 37.308f
cDVDD/287 DVDD:4069 vss 37.1817f
cDVDD/288 DVDD:4034 vss 0.413659f
cDVDD/289 DVDD:4033 vss 33.0042f
cDVDD/290 DVDD:4024 vss 0.363814f
cDVDD/291 DVDD:4014 vss 0.363814f
cDVDD/292 DVDD:4004 vss 0.363814f
cDVDD/293 DVDD:3994 vss 1.18857f
cDVDD/294 DVDD:3990 vss 0.101946f
cDVDD/295 DVDD:3986 vss 0.101946f
cDVDD/296 DVDD:3982 vss 0.101946f
cDVDD/297 DVDD:3980 vss 0.0659035f
cDVDD/298 X46/D0:neg vss 3.92581f
cDVDD/299 DVDD:2096 vss 4.85831f
cDVDD/300 DVDD:1943 vss 5.10919f
cDVDD/301 DVDD:1866 vss 4.33753f
cDVDD/302 DVDD:1787 vss 4.33755f
cDVDD/303 DVDD:1329 vss 0.810015f
cDVDD/304 DVDD:1179 vss 0.811144f
cDVDD/305 DVDD:1029 vss 0.810015f
cDVDD/306 X46/X30/D0:neg vss 10.6063f
cDVDD/307 DVDD:795 vss 7.07648f
cDVDD/308 DVDD:735 vss 4.85733f
cDVDD/309 DVDD:709 vss 0.218143f
cDVDD/310 DVDD:707 vss 4.73609f
cDVDD/311 DVDD:702 vss 7.06478f
cDVDD/312 DVDD:642 vss 0.167938f
cDVDD/313 DVDD:616 vss 0.218143f
cDVDD/314 DVDD:614 vss 0.27697f
cDVDD/315 DVDD:555 vss 3.00823f
cDVDD/316 DVDD:496 vss 2.96288f
cDVDD/317 X30/D0:neg vss 2.43325f
cDVDD/318 X29/D0:neg vss 2.50438f
cDVDD/319 X28/D0:neg vss 2.50438f
cDVDD/320 X27/D0:neg vss 2.43328f
cDVDD/321 DVDD:57 vss 3.55208f
cDVDD/322 DVDD:55 vss 3.43032f
cDVDD/323 DVDD:33 vss 0.0934477f
cDVDD/324 DVDD:31 vss 3.66223f
cDVDD/325 DVDD:28 vss 0.0936695f
cDVDD/326 DVDD:26 vss 3.4315f
cDVDD/327 DVDD:4 vss 0.0934477f
cDVDD/328 DVDD:2 vss 0.150889f
rDVDD/331 DVDD:16206 DVDD:16209 0.0113097
rDVDD/332 DVDD:16205 DVDD:16209 0.069002
rDVDD/333 DVDD:16205 DVDD:16206 0.0576923
rDVDD/334 DVDD:16200 DVDD:16206 0.0084823
rDVDD/335 DVDD:16199 DVDD:16200 0.0112876
rDVDD/336 DVDD:16195 DVDD:16200 0.0452389
rDVDD/337 DVDD:16194 DVDD:16195 0.0140333
rDVDD/338 DVDD:16176 DVDD:16177 0.00701663
rDVDD/339 DVDD:16163 DVDD 0.0118673
rDVDD/340 DVDD:16163 DVDD 0.0259005
rDVDD/341 DVDD:16157 DVDD:16160 0.0112105
rDVDD/342 DVDD:16156 DVDD:16160 0.0643601
rDVDD/343 DVDD:16156 DVDD:16157 0.0531496
rDVDD/344 DVDD:16151 DVDD:16157 0.0112105
rDVDD/345 DVDD:16150 DVDD:16151 0.0108521
rDVDD/346 DVDD:16147 DVDD:16151 0.0448421
rDVDD/347 DVDD:16146 DVDD:16147 0.0136364
rDVDD/348 DVDD:16130 DVDD:16131 0.00681818
rDVDD/349 DVDD:16117 DVDD 0.0117632
rDVDD/350 DVDD:16117 DVDD 0.0253995
rDVDD/351 DVDD:16083 DVDD:16084 0.143617
rDVDD/352 DVDD:16080 DVDD:16084 0.0365143
rDVDD/353 DVDD:16079 DVDD:16080 0.143617
rDVDD/354 DVDD:16077 DVDD:16080 0.00912857
rDVDD/355 DVDD:16076 DVDD:16079 0.00912857
rDVDD/356 DVDD:16076 DVDD:16077 0.143617
rDVDD/357 DVDD:16073 DVDD:16077 0.0456429
rDVDD/358 DVDD:16072 DVDD:16073 0.143617
rDVDD/359 DVDD:16068 DVDD:16073 0.0365143
rDVDD/360 DVDD:16067 DVDD:16072 0.0365143
rDVDD/361 DVDD:16067 DVDD:16068 0.0718085
rDVDD/362 DVDD:16065 DVDD:16068 0.0456429
rDVDD/363 DVDD:16064 DVDD:16067 0.0456429
rDVDD/364 DVDD:16064 DVDD:16065 0.143617
rDVDD/365 DVDD:16055 DVDD:16058 0.0456429
rDVDD/366 DVDD:16050 DVDD:16055 0.0456429
rDVDD/367 DVDD:16041 DVDD:16046 0.0365143
rDVDD/368 DVDD:16038 DVDD:16041 0.0456429
rDVDD/369 DVDD:16035 DVDD:16038 0.0365143
rDVDD/370 DVDD:16032 DVDD:16035 0.00912857
rDVDD/371 DVDD:16023 DVDD:16028 0.0365143
rDVDD/372 DVDD:16023 DVDD:16024 0.0718085
rDVDD/373 DVDD:16021 DVDD:16024 0.0456429
rDVDD/374 DVDD:16020 DVDD:16023 0.0456429
rDVDD/375 DVDD:16020 DVDD:16021 0.143617
rDVDD/376 DVDD:16015 DVDD:16020 0.0365143
rDVDD/377 DVDD:16006 DVDD:16011 0.0456429
rDVDD/378 DVDD:16002 DVDD:16003 0.143617
rDVDD/379 DVDD:15998 DVDD 0.0438429
rDVDD/380 DVDD:15998 DVDD:16003 0.0365143
rDVDD/381 DVDD:15997 DVDD:16002 0.0365143
rDVDD/382 DVDD:15997 DVDD:15998 0.0718085
rDVDD/383 DVDD:15990 DVDD 0.0018
rDVDD/384 DVDD:15989 DVDD 0.0018
rDVDD/385 DVDD:15989 DVDD:15990 0.143617
rDVDD/386 DVDD:15986 DVDD:15990 0.0365143
rDVDD/387 DVDD:15986 DVDD:15989 0.180131
rDVDD/388 DVDD:15976 DVDD:15977 0.143617
rDVDD/389 DVDD:15973 DVDD:15977 0.0365143
rDVDD/390 DVDD:15972 DVDD:15973 0.143617
rDVDD/391 DVDD:15970 DVDD:15973 0.00912857
rDVDD/392 DVDD:15969 DVDD:15972 0.00912857
rDVDD/393 DVDD:15969 DVDD:15970 0.143617
rDVDD/394 DVDD:15966 DVDD:15970 0.0456429
rDVDD/395 DVDD:15965 DVDD:15966 0.143617
rDVDD/396 DVDD:15961 DVDD:15966 0.0365143
rDVDD/397 DVDD:15960 DVDD:15965 0.0365143
rDVDD/398 DVDD:15960 DVDD:15961 0.0718085
rDVDD/399 DVDD:15958 DVDD:15961 0.0456429
rDVDD/400 DVDD:15957 DVDD:15960 0.0456429
rDVDD/401 DVDD:15957 DVDD:15958 0.143617
rDVDD/402 DVDD:15948 DVDD:15951 0.0456429
rDVDD/403 DVDD:15943 DVDD:15948 0.0456429
rDVDD/404 DVDD:15934 DVDD:15939 0.0365143
rDVDD/405 DVDD:15931 DVDD:15934 0.0456429
rDVDD/406 DVDD:15928 DVDD:15931 0.0365143
rDVDD/407 DVDD:15925 DVDD:15928 0.00912857
rDVDD/408 DVDD:15916 DVDD:15921 0.0365143
rDVDD/409 DVDD:15916 DVDD:15917 0.0718085
rDVDD/410 DVDD:15914 DVDD:15917 0.0456429
rDVDD/411 DVDD:15913 DVDD:15916 0.0456429
rDVDD/412 DVDD:15913 DVDD:15914 0.143617
rDVDD/413 DVDD:15908 DVDD:15913 0.0365143
rDVDD/414 DVDD:15899 DVDD:15904 0.0456429
rDVDD/415 DVDD:15895 DVDD:15896 0.143617
rDVDD/416 DVDD:15891 DVDD 0.0438429
rDVDD/417 DVDD:15891 DVDD:15896 0.0365143
rDVDD/418 DVDD:15890 DVDD:15895 0.0365143
rDVDD/419 DVDD:15890 DVDD:15891 0.0718085
rDVDD/420 DVDD:15884 DVDD 0.0018
rDVDD/421 DVDD:15883 DVDD 0.0018
rDVDD/422 DVDD:15883 DVDD:15884 0.143617
rDVDD/423 DVDD:15880 DVDD:15884 0.0365143
rDVDD/424 DVDD:15880 DVDD:15883 0.180131
rDVDD/425 DVDD:15870 DVDD:15871 0.143617
rDVDD/426 DVDD:15867 DVDD:15871 0.0365143
rDVDD/427 DVDD:15866 DVDD:15867 0.143617
rDVDD/428 DVDD:15864 DVDD:15867 0.00912857
rDVDD/429 DVDD:15863 DVDD:15866 0.00912857
rDVDD/430 DVDD:15863 DVDD:15864 0.143617
rDVDD/431 DVDD:15860 DVDD:15864 0.0456429
rDVDD/432 DVDD:15859 DVDD:15860 0.143617
rDVDD/433 DVDD:15855 DVDD:15860 0.0365143
rDVDD/434 DVDD:15854 DVDD:15859 0.0365143
rDVDD/435 DVDD:15854 DVDD:15855 0.0718085
rDVDD/436 DVDD:15852 DVDD:15855 0.0456429
rDVDD/437 DVDD:15851 DVDD:15854 0.0456429
rDVDD/438 DVDD:15851 DVDD:15852 0.143617
rDVDD/439 DVDD:15842 DVDD:15845 0.0456429
rDVDD/440 DVDD:15837 DVDD:15842 0.0456429
rDVDD/441 DVDD:15828 DVDD:15833 0.0365143
rDVDD/442 DVDD:15825 DVDD:15828 0.0456429
rDVDD/443 DVDD:15822 DVDD:15825 0.0365143
rDVDD/444 DVDD:15819 DVDD:15822 0.00912857
rDVDD/445 DVDD:15810 DVDD:15815 0.0365143
rDVDD/446 DVDD:15810 DVDD:15811 0.0718085
rDVDD/447 DVDD:15808 DVDD:15811 0.0456429
rDVDD/448 DVDD:15807 DVDD:15810 0.0456429
rDVDD/449 DVDD:15807 DVDD:15808 0.143617
rDVDD/450 DVDD:15802 DVDD:15807 0.0365143
rDVDD/451 DVDD:15793 DVDD:15798 0.0456429
rDVDD/452 DVDD:15789 DVDD:15790 0.143617
rDVDD/453 DVDD:15785 DVDD 0.0438429
rDVDD/454 DVDD:15785 DVDD:15790 0.0365143
rDVDD/455 DVDD:15784 DVDD:15789 0.0365143
rDVDD/456 DVDD:15784 DVDD:15785 0.0718085
rDVDD/457 DVDD:15777 DVDD 0.0018
rDVDD/458 DVDD:15776 DVDD 0.0018
rDVDD/459 DVDD:15776 DVDD:15777 0.143617
rDVDD/460 DVDD:15773 DVDD:15777 0.0365143
rDVDD/461 DVDD:15773 DVDD:15776 0.180131
rDVDD/462 DVDD:15741 DVDD:15749 1.5
rDVDD/463 DVDD:15740 DVDD:15741 1.5
rDVDD/464 DVDD:15737 DVDD:15743 2.25
rDVDD/465 DVDD:15737 DVDD:15741 0.0159429
rDVDD/466 DVDD:15737 DVDD:15997 0.01485
rDVDD/467 DVDD:15734 DVDD 0.00507857
rDVDD/468 DVDD:15734 DVDD:15743 1.5
rDVDD/469 DVDD:15734 DVDD:15741 0.00797143
rDVDD/470 DVDD:15733 DVDD:15737 2.25
rDVDD/471 DVDD:15733 DVDD:15734 1.5
rDVDD/472 DVDD:15724 DVDD:15729 0.0233473
rDVDD/473 DVDD:15722 DVDD:15768 0.28125
rDVDD/474 DVDD:15722 DVDD:15729 1.5
rDVDD/475 DVDD:15721 DVDD:15722 1.5
rDVDD/476 DVDD:15718 DVDD:15724 2.25
rDVDD/477 DVDD:15718 DVDD:15722 0.00489474
rDVDD/478 DVDD:15715 DVDD 0.00155921
rDVDD/479 DVDD:15715 DVDD:15724 1.5
rDVDD/480 DVDD:15715 DVDD:15722 0.00244737
rDVDD/481 DVDD:15714 DVDD:15718 2.25
rDVDD/482 DVDD:15714 DVDD:15715 1.5
rDVDD/483 DVDD:15702 DVDD:15763 0.28125
rDVDD/484 DVDD:15702 DVDD:15757 0.28125
rDVDD/485 DVDD:15702 DVDD:15753 0.28125
rDVDD/486 DVDD:15702 DVDD:15710 1.5
rDVDD/487 DVDD:15701 DVDD:15702 1.5
rDVDD/488 DVDD:15699 DVDD:15704 2.25
rDVDD/489 DVDD:15699 DVDD:15702 0.00178846
rDVDD/490 DVDD:15696 DVDD 0.000569712
rDVDD/491 DVDD:15696 DVDD:15704 1.5
rDVDD/492 DVDD:15696 DVDD:15702 0.000894231
rDVDD/493 DVDD:15695 DVDD:15701 0.0233473
rDVDD/494 DVDD:15695 DVDD:15699 2.25
rDVDD/495 DVDD:15695 DVDD:15696 1.5
rDVDD/496 DVDD:15691 DVDD:15695 0.921797
rDVDD/497 DVDD:15686 DVDD:15691 0.0233473
rDVDD/498 DVDD:15684 DVDD:15691 1.5
rDVDD/499 DVDD:15683 DVDD:15684 1.5
rDVDD/500 DVDD:15681 DVDD:15686 2.25
rDVDD/501 DVDD:15681 DVDD:15684 0.0159429
rDVDD/502 DVDD:15681 DVDD:15784 0.01485
rDVDD/503 DVDD:15678 DVDD 0.00507857
rDVDD/504 DVDD:15678 DVDD:15686 1.5
rDVDD/505 DVDD:15678 DVDD:15684 0.00797143
rDVDD/506 DVDD:15677 DVDD:15683 0.0233473
rDVDD/507 DVDD:15677 DVDD:15681 2.25
rDVDD/508 DVDD:15677 DVDD:15678 1.5
rDVDD/509 DVDD:15662 DVDD:16079 0.0225643
rDVDD/510 DVDD:15662 DVDD:15669 0.321429
rDVDD/511 DVDD:15662 DVDD:15665 0.3
rDVDD/512 DVDD:15662 DVDD:16083 0.01395
rDVDD/513 DVDD:15661 DVDD:15662 0.3
rDVDD/514 DVDD:15633 DVDD:15972 0.0225643
rDVDD/515 DVDD:15633 DVDD:15641 0.321429
rDVDD/516 DVDD:15633 DVDD:15637 0.3
rDVDD/517 DVDD:15633 DVDD:15976 0.01395
rDVDD/518 DVDD:15632 DVDD:15633 0.3
rDVDD/519 DVDD:15597 DVDD:15600 0.043937
rDVDD/520 DVDD:15591 DVDD:16199 0.00133407
rDVDD/521 DVDD:15591 DVDD:15625 0.75
rDVDD/522 DVDD:15591 DVDD:15621 0.3
rDVDD/523 DVDD:15591 DVDD:15616 0.3
rDVDD/524 DVDD:15591 DVDD:15611 0.28125
rDVDD/525 DVDD:15591 DVDD:15600 0.28125
rDVDD/526 DVDD:15591 DVDD:15597 0.75
rDVDD/527 DVDD:15591 DVDD:16205 0.00714823
rDVDD/528 DVDD:15590 DVDD:15591 0.3
rDVDD/529 DVDD:15536 DVDD:15539 0.0659055
rDVDD/530 DVDD:15534 DVDD:16150 0.004125
rDVDD/531 DVDD:15534 DVDD:15569 0.346154
rDVDD/532 DVDD:15534 DVDD:15565 0.3
rDVDD/533 DVDD:15534 DVDD:15557 0.3
rDVDD/534 DVDD:15534 DVDD:15553 0.3
rDVDD/535 DVDD:15534 DVDD:15548 0.3
rDVDD/536 DVDD:15534 DVDD:15543 0.28125
rDVDD/537 DVDD:15534 DVDD:15539 0.75
rDVDD/538 DVDD:15534 DVDD:15536 0.3
rDVDD/539 DVDD:15534 DVDD:16156 0.00708553
rDVDD/540 DVDD:15533 DVDD:15536 0.087874
rDVDD/541 DVDD:15533 DVDD:15534 0.3
rDVDD/542 DVDD:15511 DVDD:15514 0.0659055
rDVDD/543 DVDD:15484 DVDD:15487 0.0659055
rDVDD/544 DVDD:15477 DVDD:15480 0.087874
rDVDD/545 DVDD:15474 DVDD:15477 0.127559
rDVDD/546 DVDD:15471 DVDD:15474 0.043937
rDVDD/547 DVDD:15468 DVDD:15471 0.0659055
rDVDD/548 DVDD:15465 DVDD:15468 0.087874
rDVDD/549 DVDD:15462 DVDD:15465 0.0659055
rDVDD/550 DVDD:15459 DVDD:15462 0.087874
rDVDD/551 DVDD:15456 DVDD:15459 0.087874
rDVDD/552 DVDD:15453 DVDD:15456 0.127559
rDVDD/553 DVDD:15450 DVDD:15453 0.087874
rDVDD/554 DVDD:15447 DVDD:15450 0.0659055
rDVDD/555 DVDD:15444 DVDD:15447 0.087874
rDVDD/556 DVDD:15441 DVDD:15444 0.0659055
rDVDD/557 DVDD:15438 DVDD:15441 0.087874
rDVDD/558 DVDD:15436 DVDD:15523 0.346154
rDVDD/559 DVDD:15436 DVDD:15519 0.3
rDVDD/560 DVDD:15436 DVDD:15514 0.3
rDVDD/561 DVDD:15436 DVDD:15511 0.3
rDVDD/562 DVDD:15436 DVDD:15504 0.3
rDVDD/563 DVDD:15436 DVDD:15499 0.28125
rDVDD/564 DVDD:15436 DVDD:15495 0.9
rDVDD/565 DVDD:15436 DVDD:15491 0.3
rDVDD/566 DVDD:15436 DVDD:15487 0.3
rDVDD/567 DVDD:15436 DVDD:15484 0.3
rDVDD/568 DVDD:15436 DVDD:15480 0.3
rDVDD/569 DVDD:15436 DVDD:15477 0.3
rDVDD/570 DVDD:15436 DVDD:15474 0.28125
rDVDD/571 DVDD:15436 DVDD:15471 0.9
rDVDD/572 DVDD:15436 DVDD:15468 0.3
rDVDD/573 DVDD:15436 DVDD:15465 0.3
rDVDD/574 DVDD:15436 DVDD:15462 0.3
rDVDD/575 DVDD:15436 DVDD:15459 0.3
rDVDD/576 DVDD:15436 DVDD:15456 0.3
rDVDD/577 DVDD:15436 DVDD:15453 0.28125
rDVDD/578 DVDD:15436 DVDD:15450 0.346154
rDVDD/579 DVDD:15436 DVDD:15447 0.3
rDVDD/580 DVDD:15436 DVDD:15444 0.3
rDVDD/581 DVDD:15436 DVDD:15441 0.3
rDVDD/582 DVDD:15436 DVDD:15438 0.3
rDVDD/583 DVDD:15435 DVDD:15438 0.087874
rDVDD/584 DVDD:15435 DVDD:15436 0.3
rDVDD/585 DVDD:15426 DVDD:15866 0.0225643
rDVDD/586 DVDD:15426 DVDD:15435 0.54786
rDVDD/587 DVDD:15426 DVDD:15870 0.01395
rDVDD/588 DVDD:15416 DVDD:16072 0.00430714
rDVDD/589 DVDD:15416 DVDD:16076 0.0413357
rDVDD/590 DVDD:15412 DVDD:15416 1.40194
rDVDD/591 DVDD:15409 DVDD:15412 0.0659055
rDVDD/592 DVDD:15407 DVDD:15965 0.00430714
rDVDD/593 DVDD:15407 DVDD:15412 0.321429
rDVDD/594 DVDD:15407 DVDD:15409 0.3
rDVDD/595 DVDD:15407 DVDD:15969 0.0413357
rDVDD/596 DVDD:15406 DVDD:15409 0.087874
rDVDD/597 DVDD:15406 DVDD:15407 0.3
rDVDD/598 DVDD:15404 DVDD:16199 0.0188164
rDVDD/599 DVDD:15403 DVDD:15406 0.369213
rDVDD/600 DVDD:15403 DVDD:15404 2.25
rDVDD/601 DVDD:15400 DVDD:15403 0.043937
rDVDD/602 DVDD:15397 DVDD:15400 0.0659055
rDVDD/603 DVDD:15394 DVDD:15397 0.087874
rDVDD/604 DVDD:15391 DVDD:15394 0.085748
rDVDD/605 DVDD:15388 DVDD:15391 0.087874
rDVDD/606 DVDD:15385 DVDD:15388 0.0659055
rDVDD/607 DVDD:15382 DVDD:15385 0.129685
rDVDD/608 DVDD:15379 DVDD:15382 0.0659055
rDVDD/609 DVDD:15376 DVDD:15379 0.0659055
rDVDD/610 DVDD:15374 DVDD:16194 0.0239535
rDVDD/611 DVDD:15374 DVDD:15400 0.346154
rDVDD/612 DVDD:15374 DVDD:15397 0.346154
rDVDD/613 DVDD:15374 DVDD:15394 0.346154
rDVDD/614 DVDD:15374 DVDD:15391 0.346154
rDVDD/615 DVDD:15374 DVDD:15388 0.346154
rDVDD/616 DVDD:15374 DVDD:15385 0.346154
rDVDD/617 DVDD:15374 DVDD:15382 0.346154
rDVDD/618 DVDD:15374 DVDD:15379 0.346154
rDVDD/619 DVDD:15374 DVDD:15376 0.346154
rDVDD/620 DVDD:15374 DVDD:15404 0.00246903
rDVDD/621 DVDD:15373 DVDD:15376 0.0659055
rDVDD/622 DVDD:15373 DVDD:15374 0.346154
rDVDD/623 DVDD:15370 DVDD:15373 1.26248
rDVDD/624 DVDD:15367 DVDD:15370 0.0659055
rDVDD/625 DVDD:15364 DVDD:15367 0.087874
rDVDD/626 DVDD:15361 DVDD:15364 0.0659055
rDVDD/627 DVDD:15358 DVDD:15361 0.087874
rDVDD/628 DVDD:15355 DVDD:15358 0.0659055
rDVDD/629 DVDD:15352 DVDD:15355 0.087874
rDVDD/630 DVDD:15349 DVDD:15352 0.106654
rDVDD/631 DVDD:15346 DVDD:15349 0.087874
rDVDD/632 DVDD:15344 DVDD:16146 0.0265461
rDVDD/633 DVDD:15344 DVDD:15370 0.321429
rDVDD/634 DVDD:15344 DVDD:15367 0.321429
rDVDD/635 DVDD:15344 DVDD:15364 0.321429
rDVDD/636 DVDD:15344 DVDD:15361 0.321429
rDVDD/637 DVDD:15344 DVDD:15358 0.321429
rDVDD/638 DVDD:15344 DVDD:15355 0.321429
rDVDD/639 DVDD:15344 DVDD:15352 0.321429
rDVDD/640 DVDD:15344 DVDD:15349 0.321429
rDVDD/641 DVDD:15344 DVDD:15346 0.321429
rDVDD/642 DVDD:15344 DVDD:16150 0.0182961
rDVDD/643 DVDD:15343 DVDD:15346 0.0659055
rDVDD/644 DVDD:15343 DVDD:15344 0.321429
rDVDD/645 DVDD:15340 DVDD:15343 0.36815
rDVDD/646 DVDD:15337 DVDD:15340 0.0659055
rDVDD/647 DVDD:15334 DVDD:15337 0.087874
rDVDD/648 DVDD:15331 DVDD:15334 0.0659055
rDVDD/649 DVDD:15328 DVDD:15331 0.087874
rDVDD/650 DVDD:15325 DVDD:15328 0.0659055
rDVDD/651 DVDD:15322 DVDD:15325 0.087874
rDVDD/652 DVDD:15319 DVDD:15322 0.105591
rDVDD/653 DVDD:15316 DVDD:15319 0.087874
rDVDD/654 DVDD:15313 DVDD:15316 0.0659055
rDVDD/655 DVDD:15310 DVDD:15313 0.087874
rDVDD/656 DVDD:15307 DVDD:15310 0.0659055
rDVDD/657 DVDD:15304 DVDD:15307 0.087874
rDVDD/658 DVDD:15301 DVDD:15304 0.0659055
rDVDD/659 DVDD:15298 DVDD:15301 0.105591
rDVDD/660 DVDD:15295 DVDD:15298 0.087874
rDVDD/661 DVDD:15292 DVDD:15295 0.087874
rDVDD/662 DVDD:15289 DVDD:15292 0.0659055
rDVDD/663 DVDD:15286 DVDD:15289 0.087874
rDVDD/664 DVDD:15283 DVDD:15286 0.0659055
rDVDD/665 DVDD:15280 DVDD:15283 0.087874
rDVDD/666 DVDD:15277 DVDD:15280 0.083622
rDVDD/667 DVDD:15274 DVDD:15277 0.109843
rDVDD/668 DVDD:15271 DVDD:15274 0.0659055
rDVDD/669 DVDD:15268 DVDD:15271 0.087874
rDVDD/670 DVDD:15265 DVDD:15268 0.0659055
rDVDD/671 DVDD:15259 DVDD:15340 0.75
rDVDD/672 DVDD:15259 DVDD:15337 0.321429
rDVDD/673 DVDD:15259 DVDD:15334 0.321429
rDVDD/674 DVDD:15259 DVDD:15331 0.321429
rDVDD/675 DVDD:15259 DVDD:15328 0.321429
rDVDD/676 DVDD:15259 DVDD:15325 0.321429
rDVDD/677 DVDD:15259 DVDD:15322 0.321429
rDVDD/678 DVDD:15259 DVDD:15319 0.321429
rDVDD/679 DVDD:15259 DVDD:15316 0.321429
rDVDD/680 DVDD:15259 DVDD:15313 0.321429
rDVDD/681 DVDD:15259 DVDD:15310 0.321429
rDVDD/682 DVDD:15259 DVDD:15307 0.321429
rDVDD/683 DVDD:15259 DVDD:15304 0.321429
rDVDD/684 DVDD:15259 DVDD:15301 0.321429
rDVDD/685 DVDD:15259 DVDD:15298 0.321429
rDVDD/686 DVDD:15259 DVDD:15295 0.321429
rDVDD/687 DVDD:15259 DVDD:15292 0.321429
rDVDD/688 DVDD:15259 DVDD:15289 0.321429
rDVDD/689 DVDD:15259 DVDD:15286 0.321429
rDVDD/690 DVDD:15259 DVDD:15283 0.321429
rDVDD/691 DVDD:15259 DVDD:15280 0.321429
rDVDD/692 DVDD:15259 DVDD:15277 0.321429
rDVDD/693 DVDD:15259 DVDD:15274 0.321429
rDVDD/694 DVDD:15259 DVDD:15271 0.321429
rDVDD/695 DVDD:15259 DVDD:15268 0.321429
rDVDD/696 DVDD:15259 DVDD:15265 0.321429
rDVDD/697 DVDD:15259 DVDD:15261 0.321429
rDVDD/698 DVDD:15259 DVDD:15436 0.00819231
rDVDD/699 DVDD:15258 DVDD:15261 0.0659055
rDVDD/700 DVDD:15258 DVDD:15259 0.321429
rDVDD/701 DVDD:15255 DVDD:15258 0.412087
rDVDD/702 DVDD:15252 DVDD:15255 0.0659055
rDVDD/703 DVDD:15250 DVDD:15859 0.00430714
rDVDD/704 DVDD:15250 DVDD:15255 0.321429
rDVDD/705 DVDD:15250 DVDD:15252 0.3
rDVDD/706 DVDD:15250 DVDD:15863 0.0413357
rDVDD/707 DVDD:15249 DVDD:15252 0.087874
rDVDD/708 DVDD:15249 DVDD:15250 0.3
rDVDD/709 DVDD:15203 DVDD:16058 0.0134357
rDVDD/710 DVDD:15203 DVDD:15211 0.321429
rDVDD/711 DVDD:15203 DVDD:15207 0.3
rDVDD/712 DVDD:15203 DVDD:16064 0.0230786
rDVDD/713 DVDD:15202 DVDD:15203 0.3
rDVDD/714 DVDD:15174 DVDD:15951 0.0134357
rDVDD/715 DVDD:15174 DVDD:15182 0.321429
rDVDD/716 DVDD:15174 DVDD:15178 0.3
rDVDD/717 DVDD:15174 DVDD:15957 0.0230786
rDVDD/718 DVDD:15173 DVDD:15174 0.3
rDVDD/719 DVDD:15136 DVDD:15139 0.043937
rDVDD/720 DVDD:15133 DVDD:15136 0.0659055
rDVDD/721 DVDD:15129 DVDD:16188 0.0352633
rDVDD/722 DVDD:15129 DVDD:15166 0.75
rDVDD/723 DVDD:15129 DVDD:15162 0.3
rDVDD/724 DVDD:15129 DVDD:15157 0.3
rDVDD/725 DVDD:15129 DVDD:15152 0.28125
rDVDD/726 DVDD:15129 DVDD:15147 0.346154
rDVDD/727 DVDD:15129 DVDD:15143 0.3
rDVDD/728 DVDD:15129 DVDD:15139 0.28125
rDVDD/729 DVDD:15129 DVDD:15136 0.75
rDVDD/730 DVDD:15129 DVDD:15133 0.3
rDVDD/731 DVDD:15129 DVDD:16194 0.00997566
rDVDD/732 DVDD:15128 DVDD:15129 0.3
rDVDD/733 DVDD:15073 DVDD:15076 0.0659055
rDVDD/734 DVDD:15071 DVDD:16140 0.0377566
rDVDD/735 DVDD:15071 DVDD:15107 0.346154
rDVDD/736 DVDD:15071 DVDD:15103 0.3
rDVDD/737 DVDD:15071 DVDD:15098 0.3
rDVDD/738 DVDD:15071 DVDD:15094 0.3
rDVDD/739 DVDD:15071 DVDD:15090 0.3
rDVDD/740 DVDD:15071 DVDD:15085 0.3
rDVDD/741 DVDD:15071 DVDD:15080 0.28125
rDVDD/742 DVDD:15071 DVDD:15076 0.75
rDVDD/743 DVDD:15071 DVDD:15073 0.3
rDVDD/744 DVDD:15071 DVDD:16146 0.00708553
rDVDD/745 DVDD:15070 DVDD:15073 0.087874
rDVDD/746 DVDD:15070 DVDD:15071 0.3
rDVDD/747 DVDD:15048 DVDD:15051 0.0659055
rDVDD/748 DVDD:15045 DVDD:15048 0.087874
rDVDD/749 DVDD:15011 DVDD:15014 0.087874
rDVDD/750 DVDD:15004 DVDD:15007 0.043937
rDVDD/751 DVDD:15001 DVDD:15004 0.0659055
rDVDD/752 DVDD:14993 DVDD:14996 0.0659055
rDVDD/753 DVDD:14972 DVDD:14975 0.0659055
rDVDD/754 DVDD:14965 DVDD:14968 0.0659055
rDVDD/755 DVDD:14959 DVDD:15060 0.346154
rDVDD/756 DVDD:14959 DVDD:15055 0.3
rDVDD/757 DVDD:14959 DVDD:15051 0.3
rDVDD/758 DVDD:14959 DVDD:15048 0.3
rDVDD/759 DVDD:14959 DVDD:15045 0.3
rDVDD/760 DVDD:14959 DVDD:15040 0.3
rDVDD/761 DVDD:14959 DVDD:15035 0.28125
rDVDD/762 DVDD:14959 DVDD:15031 0.9
rDVDD/763 DVDD:14959 DVDD:15027 0.3
rDVDD/764 DVDD:14959 DVDD:15022 0.3
rDVDD/765 DVDD:14959 DVDD:15018 0.3
rDVDD/766 DVDD:14959 DVDD:15014 0.3
rDVDD/767 DVDD:14959 DVDD:15011 0.3
rDVDD/768 DVDD:14959 DVDD:15007 0.28125
rDVDD/769 DVDD:14959 DVDD:15004 0.9
rDVDD/770 DVDD:14959 DVDD:15001 0.3
rDVDD/771 DVDD:14959 DVDD:14996 0.3
rDVDD/772 DVDD:14959 DVDD:14993 0.3
rDVDD/773 DVDD:14959 DVDD:14988 0.3
rDVDD/774 DVDD:14959 DVDD:14984 0.3
rDVDD/775 DVDD:14959 DVDD:14980 0.28125
rDVDD/776 DVDD:14959 DVDD:14975 0.346154
rDVDD/777 DVDD:14959 DVDD:14972 0.3
rDVDD/778 DVDD:14959 DVDD:14968 0.3
rDVDD/779 DVDD:14959 DVDD:14965 0.3
rDVDD/780 DVDD:14959 DVDD:14961 0.3
rDVDD/781 DVDD:14959 DVDD:15259 0.0122885
rDVDD/782 DVDD:14958 DVDD:14961 0.087874
rDVDD/783 DVDD:14958 DVDD:14959 0.3
rDVDD/784 DVDD:14955 DVDD:14958 0.412087
rDVDD/785 DVDD:14952 DVDD:14955 0.0659055
rDVDD/786 DVDD:14950 DVDD:15845 0.0134357
rDVDD/787 DVDD:14950 DVDD:14955 0.321429
rDVDD/788 DVDD:14950 DVDD:14952 0.3
rDVDD/789 DVDD:14950 DVDD:15851 0.0230786
rDVDD/790 DVDD:14949 DVDD:14952 0.087874
rDVDD/791 DVDD:14949 DVDD:14950 0.3
rDVDD/792 DVDD:14924 DVDD:16046 0.00430714
rDVDD/793 DVDD:14924 DVDD:14932 0.321429
rDVDD/794 DVDD:14924 DVDD:14928 0.3
rDVDD/795 DVDD:14924 DVDD:16050 0.0413357
rDVDD/796 DVDD:14923 DVDD:14924 0.3
rDVDD/797 DVDD:14895 DVDD:15939 0.00430714
rDVDD/798 DVDD:14895 DVDD:14903 0.321429
rDVDD/799 DVDD:14895 DVDD:14899 0.3
rDVDD/800 DVDD:14895 DVDD:15943 0.0413357
rDVDD/801 DVDD:14894 DVDD:14895 0.3
rDVDD/802 DVDD:14888 DVDD:16188 0.00750664
rDVDD/803 DVDD:14887 DVDD:14888 2.25
rDVDD/804 DVDD:14854 DVDD:14857 0.0659055
rDVDD/805 DVDD:14847 DVDD:16183 0.0352633
rDVDD/806 DVDD:14847 DVDD:14883 0.346154
rDVDD/807 DVDD:14847 DVDD:14879 0.346154
rDVDD/808 DVDD:14847 DVDD:14874 0.346154
rDVDD/809 DVDD:14847 DVDD:14870 0.346154
rDVDD/810 DVDD:14847 DVDD:14865 0.346154
rDVDD/811 DVDD:14847 DVDD:14861 0.346154
rDVDD/812 DVDD:14847 DVDD:14857 0.346154
rDVDD/813 DVDD:14847 DVDD:14854 0.346154
rDVDD/814 DVDD:14847 DVDD:14850 0.346154
rDVDD/815 DVDD:14847 DVDD:14888 0.00246903
rDVDD/816 DVDD:14846 DVDD:14847 0.346154
rDVDD/817 DVDD:14791 DVDD:14794 0.087874
rDVDD/818 DVDD:14789 DVDD:16136 0.0377566
rDVDD/819 DVDD:14789 DVDD:14825 0.321429
rDVDD/820 DVDD:14789 DVDD:14821 0.321429
rDVDD/821 DVDD:14789 DVDD:14816 0.321429
rDVDD/822 DVDD:14789 DVDD:14812 0.321429
rDVDD/823 DVDD:14789 DVDD:14808 0.321429
rDVDD/824 DVDD:14789 DVDD:14804 0.321429
rDVDD/825 DVDD:14789 DVDD:14799 0.321429
rDVDD/826 DVDD:14789 DVDD:14794 0.321429
rDVDD/827 DVDD:14789 DVDD:14791 0.321429
rDVDD/828 DVDD:14789 DVDD:16140 0.00708553
rDVDD/829 DVDD:14788 DVDD:14791 0.0659055
rDVDD/830 DVDD:14788 DVDD:14789 0.321429
rDVDD/831 DVDD:14763 DVDD:14766 0.087874
rDVDD/832 DVDD:14729 DVDD:14732 0.087874
rDVDD/833 DVDD:14726 DVDD:14729 0.0659055
rDVDD/834 DVDD:14719 DVDD:14722 0.087874
rDVDD/835 DVDD:14711 DVDD:14714 0.0659055
rDVDD/836 DVDD:14703 DVDD:14706 0.0659055
rDVDD/837 DVDD:14695 DVDD:14698 0.083622
rDVDD/838 DVDD:14687 DVDD:14690 0.0659055
rDVDD/839 DVDD:14680 DVDD:14683 0.0659055
rDVDD/840 DVDD:14674 DVDD:16106 0.00969952
rDVDD/841 DVDD:14674 DVDD:14778 0.75
rDVDD/842 DVDD:14674 DVDD:14774 0.321429
rDVDD/843 DVDD:14674 DVDD:14770 0.321429
rDVDD/844 DVDD:14674 DVDD:14766 0.321429
rDVDD/845 DVDD:14674 DVDD:14763 0.321429
rDVDD/846 DVDD:14674 DVDD:14759 0.321429
rDVDD/847 DVDD:14674 DVDD:14754 0.321429
rDVDD/848 DVDD:14674 DVDD:14750 0.321429
rDVDD/849 DVDD:14674 DVDD:14745 0.321429
rDVDD/850 DVDD:14674 DVDD:14741 0.321429
rDVDD/851 DVDD:14674 DVDD:14736 0.321429
rDVDD/852 DVDD:14674 DVDD:14732 0.321429
rDVDD/853 DVDD:14674 DVDD:14729 0.321429
rDVDD/854 DVDD:14674 DVDD:14726 0.321429
rDVDD/855 DVDD:14674 DVDD:14722 0.321429
rDVDD/856 DVDD:14674 DVDD:14719 0.321429
rDVDD/857 DVDD:14674 DVDD:14714 0.321429
rDVDD/858 DVDD:14674 DVDD:14711 0.321429
rDVDD/859 DVDD:14674 DVDD:14706 0.321429
rDVDD/860 DVDD:14674 DVDD:14703 0.321429
rDVDD/861 DVDD:14674 DVDD:14698 0.321429
rDVDD/862 DVDD:14674 DVDD:14695 0.321429
rDVDD/863 DVDD:14674 DVDD:14690 0.321429
rDVDD/864 DVDD:14674 DVDD:14687 0.321429
rDVDD/865 DVDD:14674 DVDD:14683 0.321429
rDVDD/866 DVDD:14674 DVDD:14680 0.321429
rDVDD/867 DVDD:14674 DVDD:14676 0.321429
rDVDD/868 DVDD:14674 DVDD:14959 0.0163846
rDVDD/869 DVDD:14673 DVDD:14676 0.0659055
rDVDD/870 DVDD:14673 DVDD:14674 0.321429
rDVDD/871 DVDD:14670 DVDD:14673 0.412087
rDVDD/872 DVDD:14667 DVDD:14670 0.0659055
rDVDD/873 DVDD:14665 DVDD:15833 0.00430714
rDVDD/874 DVDD:14665 DVDD:14670 0.321429
rDVDD/875 DVDD:14665 DVDD:14667 0.3
rDVDD/876 DVDD:14665 DVDD:15837 0.0413357
rDVDD/877 DVDD:14664 DVDD:14667 0.087874
rDVDD/878 DVDD:14664 DVDD:14665 0.3
rDVDD/879 DVDD:14639 DVDD:16028 0.00572143
rDVDD/880 DVDD:14639 DVDD:14647 0.321429
rDVDD/881 DVDD:14639 DVDD:14643 0.3
rDVDD/882 DVDD:14639 DVDD:16032 0.0399214
rDVDD/883 DVDD:14638 DVDD:14639 0.3
rDVDD/884 DVDD:14610 DVDD:15921 0.00572143
rDVDD/885 DVDD:14610 DVDD:14618 0.321429
rDVDD/886 DVDD:14610 DVDD:14614 0.3
rDVDD/887 DVDD:14610 DVDD:15925 0.0399214
rDVDD/888 DVDD:14609 DVDD:14610 0.3
rDVDD/889 DVDD:14603 DVDD:16183 0.0155509
rDVDD/890 DVDD:14602 DVDD:14603 2.25
rDVDD/891 DVDD:14569 DVDD:14572 0.0659055
rDVDD/892 DVDD:14562 DVDD:16176 0.027219
rDVDD/893 DVDD:14562 DVDD:14598 0.346154
rDVDD/894 DVDD:14562 DVDD:14594 0.346154
rDVDD/895 DVDD:14562 DVDD:14589 0.346154
rDVDD/896 DVDD:14562 DVDD:14585 0.346154
rDVDD/897 DVDD:14562 DVDD:14580 0.346154
rDVDD/898 DVDD:14562 DVDD:14576 0.346154
rDVDD/899 DVDD:14562 DVDD:14572 0.346154
rDVDD/900 DVDD:14562 DVDD:14569 0.346154
rDVDD/901 DVDD:14562 DVDD:14565 0.346154
rDVDD/902 DVDD:14562 DVDD:14603 0.00246903
rDVDD/903 DVDD:14561 DVDD:14562 0.346154
rDVDD/904 DVDD:14506 DVDD:14509 0.087874
rDVDD/905 DVDD:14504 DVDD:16130 0.0297829
rDVDD/906 DVDD:14504 DVDD:14540 0.321429
rDVDD/907 DVDD:14504 DVDD:14536 0.321429
rDVDD/908 DVDD:14504 DVDD:14531 0.321429
rDVDD/909 DVDD:14504 DVDD:14527 0.321429
rDVDD/910 DVDD:14504 DVDD:14523 0.321429
rDVDD/911 DVDD:14504 DVDD:14519 0.321429
rDVDD/912 DVDD:14504 DVDD:14514 0.321429
rDVDD/913 DVDD:14504 DVDD:14509 0.321429
rDVDD/914 DVDD:14504 DVDD:14506 0.321429
rDVDD/915 DVDD:14504 DVDD:16136 0.0150592
rDVDD/916 DVDD:14503 DVDD:14506 0.0659055
rDVDD/917 DVDD:14503 DVDD:14504 0.321429
rDVDD/918 DVDD:14478 DVDD:14481 0.087874
rDVDD/919 DVDD:14444 DVDD:14447 0.087874
rDVDD/920 DVDD:14441 DVDD:14444 0.0659055
rDVDD/921 DVDD:14434 DVDD:14437 0.087874
rDVDD/922 DVDD:14426 DVDD:14429 0.0659055
rDVDD/923 DVDD:14418 DVDD:14421 0.0659055
rDVDD/924 DVDD:14410 DVDD:14413 0.083622
rDVDD/925 DVDD:14402 DVDD:14405 0.0659055
rDVDD/926 DVDD:14395 DVDD:14398 0.0659055
rDVDD/927 DVDD:14389 DVDD:14493 0.75
rDVDD/928 DVDD:14389 DVDD:14489 0.321429
rDVDD/929 DVDD:14389 DVDD:14485 0.321429
rDVDD/930 DVDD:14389 DVDD:14481 0.321429
rDVDD/931 DVDD:14389 DVDD:14478 0.321429
rDVDD/932 DVDD:14389 DVDD:14474 0.321429
rDVDD/933 DVDD:14389 DVDD:14469 0.321429
rDVDD/934 DVDD:14389 DVDD:14465 0.321429
rDVDD/935 DVDD:14389 DVDD:14460 0.321429
rDVDD/936 DVDD:14389 DVDD:14456 0.321429
rDVDD/937 DVDD:14389 DVDD:14451 0.321429
rDVDD/938 DVDD:14389 DVDD:14447 0.321429
rDVDD/939 DVDD:14389 DVDD:14444 0.321429
rDVDD/940 DVDD:14389 DVDD:14441 0.321429
rDVDD/941 DVDD:14389 DVDD:14437 0.321429
rDVDD/942 DVDD:14389 DVDD:14434 0.321429
rDVDD/943 DVDD:14389 DVDD:14429 0.321429
rDVDD/944 DVDD:14389 DVDD:14426 0.321429
rDVDD/945 DVDD:14389 DVDD:14421 0.321429
rDVDD/946 DVDD:14389 DVDD:14418 0.321429
rDVDD/947 DVDD:14389 DVDD:14413 0.321429
rDVDD/948 DVDD:14389 DVDD:14410 0.321429
rDVDD/949 DVDD:14389 DVDD:14405 0.321429
rDVDD/950 DVDD:14389 DVDD:14402 0.321429
rDVDD/951 DVDD:14389 DVDD:14398 0.321429
rDVDD/952 DVDD:14389 DVDD:14395 0.321429
rDVDD/953 DVDD:14389 DVDD:14391 0.321429
rDVDD/954 DVDD:14389 DVDD:16106 0.00959856
rDVDD/955 DVDD:14388 DVDD:14391 0.0659055
rDVDD/956 DVDD:14388 DVDD:14389 0.321429
rDVDD/957 DVDD:14385 DVDD:14388 0.412087
rDVDD/958 DVDD:14382 DVDD:14385 0.0659055
rDVDD/959 DVDD:14380 DVDD:15815 0.00572143
rDVDD/960 DVDD:14380 DVDD:14385 0.321429
rDVDD/961 DVDD:14380 DVDD:14382 0.3
rDVDD/962 DVDD:14380 DVDD:15819 0.0399214
rDVDD/963 DVDD:14379 DVDD:14382 0.087874
rDVDD/964 DVDD:14379 DVDD:14380 0.3
rDVDD/965 DVDD:14354 DVDD:16011 0.0239786
rDVDD/966 DVDD:14354 DVDD:14362 0.321429
rDVDD/967 DVDD:14354 DVDD:14358 0.3
rDVDD/968 DVDD:14354 DVDD:16015 0.0216643
rDVDD/969 DVDD:14353 DVDD:14354 0.3
rDVDD/970 DVDD:14325 DVDD:15904 0.0239786
rDVDD/971 DVDD:14325 DVDD:14333 0.321429
rDVDD/972 DVDD:14325 DVDD:14329 0.3
rDVDD/973 DVDD:14325 DVDD:15908 0.0216643
rDVDD/974 DVDD:14324 DVDD:14325 0.3
rDVDD/975 DVDD:14287 DVDD:14290 0.043937
rDVDD/976 DVDD:14284 DVDD:14287 0.0659055
rDVDD/977 DVDD:14280 DVDD:16172 0.027219
rDVDD/978 DVDD:14280 DVDD:14317 0.75
rDVDD/979 DVDD:14280 DVDD:14313 0.3
rDVDD/980 DVDD:14280 DVDD:14308 0.3
rDVDD/981 DVDD:14280 DVDD:14303 0.28125
rDVDD/982 DVDD:14280 DVDD:14298 0.346154
rDVDD/983 DVDD:14280 DVDD:14294 0.3
rDVDD/984 DVDD:14280 DVDD:14290 0.28125
rDVDD/985 DVDD:14280 DVDD:14287 0.75
rDVDD/986 DVDD:14280 DVDD:14284 0.3
rDVDD/987 DVDD:14280 DVDD:16176 0.0180199
rDVDD/988 DVDD:14279 DVDD:14280 0.3
rDVDD/989 DVDD:14224 DVDD:14227 0.0659055
rDVDD/990 DVDD:14222 DVDD:16126 0.0297829
rDVDD/991 DVDD:14222 DVDD:14258 0.346154
rDVDD/992 DVDD:14222 DVDD:14254 0.3
rDVDD/993 DVDD:14222 DVDD:14249 0.3
rDVDD/994 DVDD:14222 DVDD:14245 0.3
rDVDD/995 DVDD:14222 DVDD:14241 0.3
rDVDD/996 DVDD:14222 DVDD:14236 0.3
rDVDD/997 DVDD:14222 DVDD:14231 0.28125
rDVDD/998 DVDD:14222 DVDD:14227 0.75
rDVDD/999 DVDD:14222 DVDD:14224 0.3
rDVDD/1000 DVDD:14222 DVDD:16130 0.0150592
rDVDD/1001 DVDD:14221 DVDD:14224 0.087874
rDVDD/1002 DVDD:14221 DVDD:14222 0.3
rDVDD/1003 DVDD:14199 DVDD:14202 0.0659055
rDVDD/1004 DVDD:14196 DVDD:14199 0.087874
rDVDD/1005 DVDD:14162 DVDD:14165 0.087874
rDVDD/1006 DVDD:14155 DVDD:14158 0.043937
rDVDD/1007 DVDD:14152 DVDD:14155 0.0659055
rDVDD/1008 DVDD:14144 DVDD:14147 0.0659055
rDVDD/1009 DVDD:14123 DVDD:14126 0.0659055
rDVDD/1010 DVDD:14116 DVDD:14119 0.0659055
rDVDD/1011 DVDD:14110 DVDD:14211 0.346154
rDVDD/1012 DVDD:14110 DVDD:14206 0.3
rDVDD/1013 DVDD:14110 DVDD:14202 0.3
rDVDD/1014 DVDD:14110 DVDD:14199 0.3
rDVDD/1015 DVDD:14110 DVDD:14196 0.3
rDVDD/1016 DVDD:14110 DVDD:14191 0.3
rDVDD/1017 DVDD:14110 DVDD:14186 0.28125
rDVDD/1018 DVDD:14110 DVDD:14182 0.9
rDVDD/1019 DVDD:14110 DVDD:14178 0.3
rDVDD/1020 DVDD:14110 DVDD:14173 0.3
rDVDD/1021 DVDD:14110 DVDD:14169 0.3
rDVDD/1022 DVDD:14110 DVDD:14165 0.3
rDVDD/1023 DVDD:14110 DVDD:14162 0.3
rDVDD/1024 DVDD:14110 DVDD:14158 0.28125
rDVDD/1025 DVDD:14110 DVDD:14155 0.9
rDVDD/1026 DVDD:14110 DVDD:14152 0.3
rDVDD/1027 DVDD:14110 DVDD:14147 0.3
rDVDD/1028 DVDD:14110 DVDD:14144 0.3
rDVDD/1029 DVDD:14110 DVDD:14139 0.3
rDVDD/1030 DVDD:14110 DVDD:14135 0.3
rDVDD/1031 DVDD:14110 DVDD:14131 0.28125
rDVDD/1032 DVDD:14110 DVDD:14126 0.346154
rDVDD/1033 DVDD:14110 DVDD:14123 0.3
rDVDD/1034 DVDD:14110 DVDD:14119 0.3
rDVDD/1035 DVDD:14110 DVDD:14116 0.3
rDVDD/1036 DVDD:14110 DVDD:14112 0.3
rDVDD/1037 DVDD:14110 DVDD:14389 0.0163846
rDVDD/1038 DVDD:14109 DVDD:14112 0.087874
rDVDD/1039 DVDD:14109 DVDD:14110 0.3
rDVDD/1040 DVDD:14106 DVDD:14109 0.412087
rDVDD/1041 DVDD:14103 DVDD:14106 0.0659055
rDVDD/1042 DVDD:14101 DVDD:15798 0.0239786
rDVDD/1043 DVDD:14101 DVDD:14106 0.321429
rDVDD/1044 DVDD:14101 DVDD:14103 0.3
rDVDD/1045 DVDD:14101 DVDD:15802 0.0216643
rDVDD/1046 DVDD:14100 DVDD:14103 0.087874
rDVDD/1047 DVDD:14100 DVDD:14101 0.3
rDVDD/1048 DVDD:14082 DVDD:16002 0.00572143
rDVDD/1049 DVDD:14082 DVDD:16006 0.0399214
rDVDD/1050 DVDD:14078 DVDD:14082 1.40194
rDVDD/1051 DVDD:14075 DVDD:14078 0.0659055
rDVDD/1052 DVDD:14073 DVDD:15895 0.00572143
rDVDD/1053 DVDD:14073 DVDD:14078 0.321429
rDVDD/1054 DVDD:14073 DVDD:14075 0.3
rDVDD/1055 DVDD:14073 DVDD:15899 0.0399214
rDVDD/1056 DVDD:14072 DVDD:14075 0.087874
rDVDD/1057 DVDD:14072 DVDD:14073 0.3
rDVDD/1058 DVDD:14070 DVDD:16172 0.00424115
rDVDD/1059 DVDD:14069 DVDD:14072 0.369213
rDVDD/1060 DVDD:14069 DVDD:14070 2.25
rDVDD/1061 DVDD:14066 DVDD:14069 0.043937
rDVDD/1062 DVDD:14063 DVDD:14066 0.0659055
rDVDD/1063 DVDD:14060 DVDD:14063 0.087874
rDVDD/1064 DVDD:14057 DVDD:14060 0.085748
rDVDD/1065 DVDD:14054 DVDD:14057 0.087874
rDVDD/1066 DVDD:14051 DVDD:14054 0.0659055
rDVDD/1067 DVDD:14048 DVDD:14051 0.129685
rDVDD/1068 DVDD:14045 DVDD:14048 0.0659055
rDVDD/1069 DVDD:14042 DVDD:14045 0.0659055
rDVDD/1070 DVDD:14040 DVDD:14066 0.346154
rDVDD/1071 DVDD:14040 DVDD:14063 0.346154
rDVDD/1072 DVDD:14040 DVDD:14060 0.346154
rDVDD/1073 DVDD:14040 DVDD:14057 0.346154
rDVDD/1074 DVDD:14040 DVDD:14054 0.346154
rDVDD/1075 DVDD:14040 DVDD:14051 0.346154
rDVDD/1076 DVDD:14040 DVDD:14048 0.346154
rDVDD/1077 DVDD:14040 DVDD:14045 0.346154
rDVDD/1078 DVDD:14040 DVDD:14042 0.346154
rDVDD/1079 DVDD:14040 DVDD:14070 0.00246903
rDVDD/1080 DVDD:14039 DVDD:14042 0.0659055
rDVDD/1081 DVDD:14039 DVDD:14040 0.346154
rDVDD/1082 DVDD:14036 DVDD:14039 1.26248
rDVDD/1083 DVDD:14033 DVDD:14036 0.0659055
rDVDD/1084 DVDD:14030 DVDD:14033 0.087874
rDVDD/1085 DVDD:14027 DVDD:14030 0.0659055
rDVDD/1086 DVDD:14024 DVDD:14027 0.087874
rDVDD/1087 DVDD:14021 DVDD:14024 0.0659055
rDVDD/1088 DVDD:14018 DVDD:14021 0.087874
rDVDD/1089 DVDD:14015 DVDD:14018 0.106654
rDVDD/1090 DVDD:14012 DVDD:14015 0.087874
rDVDD/1091 DVDD:14010 DVDD:15718 0.0175263
rDVDD/1092 DVDD:14010 DVDD:14036 0.321429
rDVDD/1093 DVDD:14010 DVDD:14033 0.321429
rDVDD/1094 DVDD:14010 DVDD:14030 0.321429
rDVDD/1095 DVDD:14010 DVDD:14027 0.321429
rDVDD/1096 DVDD:14010 DVDD:14024 0.321429
rDVDD/1097 DVDD:14010 DVDD:14021 0.321429
rDVDD/1098 DVDD:14010 DVDD:14018 0.321429
rDVDD/1099 DVDD:14010 DVDD:14015 0.321429
rDVDD/1100 DVDD:14010 DVDD:14012 0.321429
rDVDD/1101 DVDD:14010 DVDD:16126 0.00384868
rDVDD/1102 DVDD:14009 DVDD:14012 0.0659055
rDVDD/1103 DVDD:14009 DVDD:14010 0.321429
rDVDD/1104 DVDD:14006 DVDD:14009 0.36815
rDVDD/1105 DVDD:14003 DVDD:14006 0.0659055
rDVDD/1106 DVDD:14000 DVDD:14003 0.087874
rDVDD/1107 DVDD:13997 DVDD:14000 0.0659055
rDVDD/1108 DVDD:13994 DVDD:13997 0.087874
rDVDD/1109 DVDD:13991 DVDD:13994 0.0659055
rDVDD/1110 DVDD:13988 DVDD:13991 0.087874
rDVDD/1111 DVDD:13985 DVDD:13988 0.105591
rDVDD/1112 DVDD:13982 DVDD:13985 0.087874
rDVDD/1113 DVDD:13979 DVDD:13982 0.0659055
rDVDD/1114 DVDD:13976 DVDD:13979 0.087874
rDVDD/1115 DVDD:13973 DVDD:13976 0.0659055
rDVDD/1116 DVDD:13970 DVDD:13973 0.087874
rDVDD/1117 DVDD:13967 DVDD:13970 0.0659055
rDVDD/1118 DVDD:13964 DVDD:13967 0.105591
rDVDD/1119 DVDD:13961 DVDD:13964 0.087874
rDVDD/1120 DVDD:13958 DVDD:13961 0.087874
rDVDD/1121 DVDD:13955 DVDD:13958 0.0659055
rDVDD/1122 DVDD:13952 DVDD:13955 0.087874
rDVDD/1123 DVDD:13949 DVDD:13952 0.0659055
rDVDD/1124 DVDD:13946 DVDD:13949 0.087874
rDVDD/1125 DVDD:13943 DVDD:13946 0.083622
rDVDD/1126 DVDD:13940 DVDD:13943 0.109843
rDVDD/1127 DVDD:13937 DVDD:13940 0.0659055
rDVDD/1128 DVDD:13934 DVDD:13937 0.087874
rDVDD/1129 DVDD:13931 DVDD:13934 0.0659055
rDVDD/1130 DVDD:13925 DVDD:15699 0.00640385
rDVDD/1131 DVDD:13925 DVDD:14006 0.75
rDVDD/1132 DVDD:13925 DVDD:14003 0.321429
rDVDD/1133 DVDD:13925 DVDD:14000 0.321429
rDVDD/1134 DVDD:13925 DVDD:13997 0.321429
rDVDD/1135 DVDD:13925 DVDD:13994 0.321429
rDVDD/1136 DVDD:13925 DVDD:13991 0.321429
rDVDD/1137 DVDD:13925 DVDD:13988 0.321429
rDVDD/1138 DVDD:13925 DVDD:13985 0.321429
rDVDD/1139 DVDD:13925 DVDD:13982 0.321429
rDVDD/1140 DVDD:13925 DVDD:13979 0.321429
rDVDD/1141 DVDD:13925 DVDD:13976 0.321429
rDVDD/1142 DVDD:13925 DVDD:13973 0.321429
rDVDD/1143 DVDD:13925 DVDD:13970 0.321429
rDVDD/1144 DVDD:13925 DVDD:13967 0.321429
rDVDD/1145 DVDD:13925 DVDD:13964 0.321429
rDVDD/1146 DVDD:13925 DVDD:13961 0.321429
rDVDD/1147 DVDD:13925 DVDD:13958 0.321429
rDVDD/1148 DVDD:13925 DVDD:13955 0.321429
rDVDD/1149 DVDD:13925 DVDD:13952 0.321429
rDVDD/1150 DVDD:13925 DVDD:13949 0.321429
rDVDD/1151 DVDD:13925 DVDD:13946 0.321429
rDVDD/1152 DVDD:13925 DVDD:13943 0.321429
rDVDD/1153 DVDD:13925 DVDD:13940 0.321429
rDVDD/1154 DVDD:13925 DVDD:13937 0.321429
rDVDD/1155 DVDD:13925 DVDD:13934 0.321429
rDVDD/1156 DVDD:13925 DVDD:13931 0.321429
rDVDD/1157 DVDD:13925 DVDD:13927 0.321429
rDVDD/1158 DVDD:13925 DVDD:14110 0.0122885
rDVDD/1159 DVDD:13924 DVDD:13927 0.0659055
rDVDD/1160 DVDD:13924 DVDD:13925 0.321429
rDVDD/1161 DVDD:13921 DVDD:13924 0.412087
rDVDD/1162 DVDD:13918 DVDD:13921 0.0659055
rDVDD/1163 DVDD:13916 DVDD:15789 0.00572143
rDVDD/1164 DVDD:13916 DVDD:13921 0.321429
rDVDD/1165 DVDD:13916 DVDD:13918 0.3
rDVDD/1166 DVDD:13916 DVDD:15793 0.0399214
rDVDD/1167 DVDD:13915 DVDD:13918 0.087874
rDVDD/1168 DVDD:13915 DVDD:13916 0.3
rDVDD/1169 DVDD:13859 DVDD:15890 0.0129214
rDVDD/1170 DVDD:13858 DVDD:13859 4.5
rDVDD/1171 DVDD:13834 DVDD 0.02295
rDVDD/1172 DVDD:13834 DVDD:13854 1.5
rDVDD/1173 DVDD:13834 DVDD:13847 1.5
rDVDD/1174 DVDD:13834 DVDD:13840 1.5
rDVDD/1175 DVDD:13834 DVDD:13859 0.00797143
rDVDD/1176 DVDD:13833 DVDD:13834 1.5
rDVDD/1177 DVDD:13770 DVDD:13773 0.0558
rDVDD/1178 DVDD:13767 DVDD:13770 0.1116
rDVDD/1179 DVDD:13753 DVDD 0.00710841
rDVDD/1180 DVDD:13753 DVDD:13800 1.5
rDVDD/1181 DVDD:13753 DVDD:13793 1.5
rDVDD/1182 DVDD:13753 DVDD:13786 1.5
rDVDD/1183 DVDD:13753 DVDD:13779 1.5
rDVDD/1184 DVDD:13753 DVDD:13773 1.5
rDVDD/1185 DVDD:13753 DVDD:13770 1.5
rDVDD/1186 DVDD:13753 DVDD:13767 1.5
rDVDD/1187 DVDD:13753 DVDD:13759 1.5
rDVDD/1188 DVDD:13753 DVDD:14040 0.0195531
rDVDD/1189 DVDD:13752 DVDD:13753 1.5
rDVDD/1190 DVDD:13735 DVDD:15741 0.346154
rDVDD/1191 DVDD:13731 DVDD:15741 0.3
rDVDD/1192 DVDD:13725 DVDD:15724 0.0233473
rDVDD/1193 DVDD:13725 DVDD:15722 0.9
rDVDD/1194 DVDD:13720 DVDD:15722 0.3
rDVDD/1195 DVDD:13716 DVDD:15722 0.3
rDVDD/1196 DVDD:13712 DVDD:15722 0.3
rDVDD/1197 DVDD:13707 DVDD:15722 0.3
rDVDD/1198 DVDD:13703 DVDD:15722 0.3
rDVDD/1199 DVDD:13698 DVDD:15722 0.346154
rDVDD/1200 DVDD:13695 DVDD:15721 0.0466946
rDVDD/1201 DVDD:13695 DVDD:13698 0.0700418
rDVDD/1202 DVDD:13695 DVDD:15722 0.3
rDVDD/1203 DVDD:13690 DVDD:15704 0.0233473
rDVDD/1204 DVDD:13690 DVDD:15702 0.9
rDVDD/1205 DVDD:13686 DVDD:15702 0.3
rDVDD/1206 DVDD:13681 DVDD:15702 0.3
rDVDD/1207 DVDD:13678 DVDD:13681 0.0700418
rDVDD/1208 DVDD:13678 DVDD:15702 0.3
rDVDD/1209 DVDD:13675 DVDD:13678 0.0933891
rDVDD/1210 DVDD:13675 DVDD:15702 0.3
rDVDD/1211 DVDD:13670 DVDD:15702 0.3
rDVDD/1212 DVDD:13665 DVDD:15702 0.9
rDVDD/1213 DVDD:13661 DVDD:15702 0.3
rDVDD/1214 DVDD:13656 DVDD:15702 0.3
rDVDD/1215 DVDD:13652 DVDD:15702 0.3
rDVDD/1216 DVDD:13648 DVDD:15702 0.3
rDVDD/1217 DVDD:13645 DVDD:13648 0.0933891
rDVDD/1218 DVDD:13645 DVDD:15702 0.3
rDVDD/1219 DVDD:13645 DVDD:15757 0.269139
rDVDD/1220 DVDD:13641 DVDD:15757 0.0466946
rDVDD/1221 DVDD:13641 DVDD:15702 0.9
rDVDD/1222 DVDD:13638 DVDD:13641 0.0700418
rDVDD/1223 DVDD:13638 DVDD:15702 0.3
rDVDD/1224 DVDD:13635 DVDD:13638 0.0933891
rDVDD/1225 DVDD:13635 DVDD:15702 0.3
rDVDD/1226 DVDD:13632 DVDD:13635 0.0700418
rDVDD/1227 DVDD:13632 DVDD:15702 0.3
rDVDD/1228 DVDD:13629 DVDD:13632 0.0933891
rDVDD/1229 DVDD:13629 DVDD:15702 0.3
rDVDD/1230 DVDD:13626 DVDD:13629 0.0933891
rDVDD/1231 DVDD:13626 DVDD:15702 0.3
rDVDD/1232 DVDD:13626 DVDD:15753 0.269139
rDVDD/1233 DVDD:13622 DVDD:15753 0.0466946
rDVDD/1234 DVDD:13622 DVDD:15702 0.9
rDVDD/1235 DVDD:13619 DVDD:13622 0.0700418
rDVDD/1236 DVDD:13619 DVDD:15702 0.3
rDVDD/1237 DVDD:13616 DVDD:13619 0.0933891
rDVDD/1238 DVDD:13616 DVDD:15702 0.3
rDVDD/1239 DVDD:13613 DVDD:13616 0.0700418
rDVDD/1240 DVDD:13613 DVDD:15702 0.3
rDVDD/1241 DVDD:13610 DVDD:13613 0.0933891
rDVDD/1242 DVDD:13610 DVDD:15702 0.3
rDVDD/1243 DVDD:13607 DVDD:15701 0.0466946
rDVDD/1244 DVDD:13607 DVDD:13610 0.0933891
rDVDD/1245 DVDD:13607 DVDD:15702 0.3
rDVDD/1246 DVDD:13602 DVDD:15686 0.0700418
rDVDD/1247 DVDD:13602 DVDD:15684 0.346154
rDVDD/1248 DVDD:13599 DVDD:15683 0.0466946
rDVDD/1249 DVDD:13599 DVDD:13602 0.0700418
rDVDD/1250 DVDD:13599 DVDD:15684 0.3
rDVDD/1251 DVDD:13590 DVDD:13592 0.793937
rDVDD/1252 DVDD:13589 DVDD:13592 0.02232
rDVDD/1253 DVDD:13589 DVDD:13590 0.5625
rDVDD/1254 DVDD:13587 DVDD:13590 0.0659055
rDVDD/1255 DVDD:13586 DVDD:13589 0.03348
rDVDD/1256 DVDD:13586 DVDD:13587 0.5625
rDVDD/1257 DVDD:13584 DVDD:15669 0.0242717
rDVDD/1258 DVDD:13584 DVDD:13587 0.043937
rDVDD/1259 DVDD:13583 DVDD:13586 0.02232
rDVDD/1260 DVDD:13583 DVDD:13584 0.5625
rDVDD/1261 DVDD:13581 DVDD:15665 0.0242717
rDVDD/1262 DVDD:13581 DVDD:15669 0.0416339
rDVDD/1263 DVDD:13580 DVDD:13583 0.03348
rDVDD/1264 DVDD:13580 DVDD:13581 0.5625
rDVDD/1265 DVDD:13578 DVDD:15661 0.0462402
rDVDD/1266 DVDD:13578 DVDD:15665 0.0416339
rDVDD/1267 DVDD:13577 DVDD:13580 0.03348
rDVDD/1268 DVDD:13577 DVDD:13578 0.5625
rDVDD/1269 DVDD:13574 DVDD:13577 0.02232
rDVDD/1270 DVDD:13574 DVDD:15661 0.5625
rDVDD/1271 DVDD:13572 DVDD:15661 0.0636024
rDVDD/1272 DVDD:13571 DVDD:13574 0.03348
rDVDD/1273 DVDD:13571 DVDD:13572 0.5625
rDVDD/1274 DVDD:13569 DVDD:13572 0.0659055
rDVDD/1275 DVDD:13568 DVDD:13571 0.03348
rDVDD/1276 DVDD:13568 DVDD:13569 0.5625
rDVDD/1277 DVDD:13566 DVDD:13569 0.043937
rDVDD/1278 DVDD:13565 DVDD:13568 0.02232
rDVDD/1279 DVDD:13565 DVDD:13566 0.5625
rDVDD/1280 DVDD:13558 DVDD:13566 0.194173
rDVDD/1281 DVDD:13557 DVDD:13558 0.75
rDVDD/1282 DVDD:13555 DVDD:13558 0.043937
rDVDD/1283 DVDD:13554 DVDD:13557 0.02232
rDVDD/1284 DVDD:13554 DVDD:13555 0.5625
rDVDD/1285 DVDD:13552 DVDD:13555 0.0659055
rDVDD/1286 DVDD:13551 DVDD:13554 0.03348
rDVDD/1287 DVDD:13551 DVDD:13552 0.5625
rDVDD/1288 DVDD:13549 DVDD:13552 0.043937
rDVDD/1289 DVDD:13548 DVDD:13551 0.02232
rDVDD/1290 DVDD:13548 DVDD:13549 0.5625
rDVDD/1291 DVDD:13546 DVDD:13549 0.0659055
rDVDD/1292 DVDD:13545 DVDD:13548 0.03348
rDVDD/1293 DVDD:13545 DVDD:13546 0.5625
rDVDD/1294 DVDD:13543 DVDD:13546 0.0659055
rDVDD/1295 DVDD:13542 DVDD:13545 0.03348
rDVDD/1296 DVDD:13542 DVDD:13543 0.5625
rDVDD/1297 DVDD:13540 DVDD:13543 0.043937
rDVDD/1298 DVDD:13539 DVDD:13542 0.02232
rDVDD/1299 DVDD:13539 DVDD:13540 0.5625
rDVDD/1300 DVDD:13537 DVDD:13540 0.0659055
rDVDD/1301 DVDD:13536 DVDD:13539 0.03348
rDVDD/1302 DVDD:13536 DVDD:13537 0.5625
rDVDD/1303 DVDD:13534 DVDD:13537 0.0659055
rDVDD/1304 DVDD:13533 DVDD:13536 0.03348
rDVDD/1305 DVDD:13533 DVDD:13534 0.5625
rDVDD/1306 DVDD:13531 DVDD:13534 0.043937
rDVDD/1307 DVDD:13530 DVDD:13533 0.02232
rDVDD/1308 DVDD:13530 DVDD:13531 0.5625
rDVDD/1309 DVDD:13523 DVDD:13531 0.194173
rDVDD/1310 DVDD:13522 DVDD:13523 0.75
rDVDD/1311 DVDD:13520 DVDD:13523 0.043937
rDVDD/1312 DVDD:13519 DVDD:13522 0.02232
rDVDD/1313 DVDD:13519 DVDD:13520 0.5625
rDVDD/1314 DVDD:13517 DVDD:13520 0.0659055
rDVDD/1315 DVDD:13516 DVDD:13519 0.03348
rDVDD/1316 DVDD:13516 DVDD:13517 0.5625
rDVDD/1317 DVDD:13514 DVDD:15641 0.0426969
rDVDD/1318 DVDD:13514 DVDD:13517 0.043937
rDVDD/1319 DVDD:13513 DVDD:13516 0.02232
rDVDD/1320 DVDD:13513 DVDD:13514 0.5625
rDVDD/1321 DVDD:13511 DVDD:15637 0.0426969
rDVDD/1322 DVDD:13511 DVDD:15641 0.0232087
rDVDD/1323 DVDD:13510 DVDD:13513 0.03348
rDVDD/1324 DVDD:13510 DVDD:13511 0.5625
rDVDD/1325 DVDD:13508 DVDD:15637 0.0232087
rDVDD/1326 DVDD:13507 DVDD:13510 0.03348
rDVDD/1327 DVDD:13507 DVDD:13508 0.5625
rDVDD/1328 DVDD:13505 DVDD:15632 0.0207283
rDVDD/1329 DVDD:13505 DVDD:13508 0.043937
rDVDD/1330 DVDD:13504 DVDD:13507 0.02232
rDVDD/1331 DVDD:13504 DVDD:13505 0.5625
rDVDD/1332 DVDD:13502 DVDD:15632 0.0451772
rDVDD/1333 DVDD:13501 DVDD:13504 0.03348
rDVDD/1334 DVDD:13501 DVDD:13502 0.5625
rDVDD/1335 DVDD:13499 DVDD:13502 0.0659055
rDVDD/1336 DVDD:13498 DVDD:13501 0.03348
rDVDD/1337 DVDD:13498 DVDD:13499 0.5625
rDVDD/1338 DVDD:13496 DVDD:13499 0.043937
rDVDD/1339 DVDD:13495 DVDD:13498 0.02232
rDVDD/1340 DVDD:13495 DVDD:13496 0.5625
rDVDD/1341 DVDD:13488 DVDD:15625 0.0200197
rDVDD/1342 DVDD:13488 DVDD:13496 0.194173
rDVDD/1343 DVDD:13487 DVDD:13488 0.75
rDVDD/1344 DVDD:13485 DVDD:15621 0.0419882
rDVDD/1345 DVDD:13485 DVDD:15625 0.0239173
rDVDD/1346 DVDD:13484 DVDD:13487 0.02232
rDVDD/1347 DVDD:13484 DVDD:13485 0.5625
rDVDD/1348 DVDD:13482 DVDD:15621 0.0239173
rDVDD/1349 DVDD:13481 DVDD:13484 0.03348
rDVDD/1350 DVDD:13481 DVDD:13482 0.5625
rDVDD/1351 DVDD:13479 DVDD:15616 0.0200197
rDVDD/1352 DVDD:13479 DVDD:13482 0.043937
rDVDD/1353 DVDD:13478 DVDD:13481 0.02232
rDVDD/1354 DVDD:13478 DVDD:13479 0.5625
rDVDD/1355 DVDD:13476 DVDD:15616 0.0458858
rDVDD/1356 DVDD:13475 DVDD:13478 0.03348
rDVDD/1357 DVDD:13475 DVDD:13476 0.5625
rDVDD/1358 DVDD:13473 DVDD:15611 0.0178937
rDVDD/1359 DVDD:13473 DVDD:13476 0.0659055
rDVDD/1360 DVDD:13472 DVDD:13475 0.03348
rDVDD/1361 DVDD:13472 DVDD:13473 0.5625
rDVDD/1362 DVDD:13470 DVDD:15611 0.0260433
rDVDD/1363 DVDD:13469 DVDD:13472 0.02232
rDVDD/1364 DVDD:13469 DVDD:13470 0.5625
rDVDD/1365 DVDD:13467 DVDD:13470 0.0659055
rDVDD/1366 DVDD:13467 DVDD:15591 0.346154
rDVDD/1367 DVDD:13466 DVDD:13469 0.03348
rDVDD/1368 DVDD:13466 DVDD:13467 0.5625
rDVDD/1369 DVDD:13464 DVDD:13467 0.0659055
rDVDD/1370 DVDD:13464 DVDD:15591 0.3
rDVDD/1371 DVDD:13463 DVDD:13466 0.03348
rDVDD/1372 DVDD:13463 DVDD:13464 0.5625
rDVDD/1373 DVDD:13461 DVDD:15600 0.0816732
rDVDD/1374 DVDD:13461 DVDD:13464 0.043937
rDVDD/1375 DVDD:13460 DVDD:13463 0.02232
rDVDD/1376 DVDD:13460 DVDD:13461 0.5625
rDVDD/1377 DVDD:13453 DVDD:15597 0.068563
rDVDD/1378 DVDD:13453 DVDD:15591 0.3
rDVDD/1379 DVDD:13452 DVDD:13453 0.75
rDVDD/1380 DVDD:13450 DVDD:15590 0.0412795
rDVDD/1381 DVDD:13450 DVDD:13453 0.043937
rDVDD/1382 DVDD:13449 DVDD:13452 0.02232
rDVDD/1383 DVDD:13449 DVDD:13450 0.5625
rDVDD/1384 DVDD:13447 DVDD:15590 0.024626
rDVDD/1385 DVDD:13446 DVDD:13449 0.03348
rDVDD/1386 DVDD:13446 DVDD:13447 0.5625
rDVDD/1387 DVDD:13444 DVDD:13447 0.043937
rDVDD/1388 DVDD:13443 DVDD:13446 0.02232
rDVDD/1389 DVDD:13443 DVDD:13444 0.5625
rDVDD/1390 DVDD:13441 DVDD:13444 0.0659055
rDVDD/1391 DVDD:13440 DVDD:13443 0.03348
rDVDD/1392 DVDD:13440 DVDD:13441 0.5625
rDVDD/1393 DVDD:13438 DVDD:13441 0.0659055
rDVDD/1394 DVDD:13437 DVDD:13440 0.03348
rDVDD/1395 DVDD:13437 DVDD:13438 0.5625
rDVDD/1396 DVDD:13435 DVDD:13438 0.043937
rDVDD/1397 DVDD:13434 DVDD:13437 0.02232
rDVDD/1398 DVDD:13434 DVDD:13435 0.5625
rDVDD/1399 DVDD:13432 DVDD:13435 0.0659055
rDVDD/1400 DVDD:13431 DVDD:13434 0.03348
rDVDD/1401 DVDD:13431 DVDD:13432 0.5625
rDVDD/1402 DVDD:13429 DVDD:13432 0.0659055
rDVDD/1403 DVDD:13428 DVDD:13431 0.03348
rDVDD/1404 DVDD:13428 DVDD:13429 0.5625
rDVDD/1405 DVDD:13426 DVDD:13429 0.043937
rDVDD/1406 DVDD:13425 DVDD:13428 0.02232
rDVDD/1407 DVDD:13425 DVDD:13426 0.5625
rDVDD/1408 DVDD:13418 DVDD:13426 0.194173
rDVDD/1409 DVDD:13417 DVDD:13418 0.75
rDVDD/1410 DVDD:13415 DVDD:13418 0.043937
rDVDD/1411 DVDD:13414 DVDD:13417 0.02232
rDVDD/1412 DVDD:13414 DVDD:13415 0.5625
rDVDD/1413 DVDD:13412 DVDD:13415 0.0659055
rDVDD/1414 DVDD:13411 DVDD:13414 0.03348
rDVDD/1415 DVDD:13411 DVDD:13412 0.5625
rDVDD/1416 DVDD:13409 DVDD:13412 0.043937
rDVDD/1417 DVDD:13408 DVDD:13411 0.02232
rDVDD/1418 DVDD:13408 DVDD:13409 0.5625
rDVDD/1419 DVDD:13406 DVDD:13409 0.0659055
rDVDD/1420 DVDD:13405 DVDD:13408 0.03348
rDVDD/1421 DVDD:13405 DVDD:13406 0.5625
rDVDD/1422 DVDD:13403 DVDD:13406 0.0659055
rDVDD/1423 DVDD:13402 DVDD:13405 0.03348
rDVDD/1424 DVDD:13402 DVDD:13403 0.5625
rDVDD/1425 DVDD:13400 DVDD:13403 0.043937
rDVDD/1426 DVDD:13399 DVDD:13402 0.02232
rDVDD/1427 DVDD:13399 DVDD:13400 0.5625
rDVDD/1428 DVDD:13397 DVDD:13400 0.0659055
rDVDD/1429 DVDD:13396 DVDD:13399 0.03348
rDVDD/1430 DVDD:13396 DVDD:13397 0.5625
rDVDD/1431 DVDD:13394 DVDD:13397 0.0659055
rDVDD/1432 DVDD:13393 DVDD:13396 0.03348
rDVDD/1433 DVDD:13393 DVDD:13394 0.5625
rDVDD/1434 DVDD:13391 DVDD:15569 0.142972
rDVDD/1435 DVDD:13391 DVDD:13394 0.043937
rDVDD/1436 DVDD:13390 DVDD:13393 0.02232
rDVDD/1437 DVDD:13390 DVDD:13391 0.5625
rDVDD/1438 DVDD:13383 DVDD:15565 0.0147047
rDVDD/1439 DVDD:13383 DVDD:15569 0.0512008
rDVDD/1440 DVDD:13382 DVDD:13383 0.75
rDVDD/1441 DVDD:13380 DVDD:15565 0.0292323
rDVDD/1442 DVDD:13379 DVDD:13382 0.02232
rDVDD/1443 DVDD:13379 DVDD:13380 0.5625
rDVDD/1444 DVDD:13377 DVDD:13380 0.0659055
rDVDD/1445 DVDD:13377 DVDD:15534 0.3
rDVDD/1446 DVDD:13376 DVDD:13379 0.03348
rDVDD/1447 DVDD:13376 DVDD:13377 0.5625
rDVDD/1448 DVDD:13374 DVDD:15557 0.0147047
rDVDD/1449 DVDD:13374 DVDD:13377 0.043937
rDVDD/1450 DVDD:13373 DVDD:13376 0.02232
rDVDD/1451 DVDD:13373 DVDD:13374 0.5625
rDVDD/1452 DVDD:13371 DVDD:15553 0.0366732
rDVDD/1453 DVDD:13371 DVDD:15557 0.0512008
rDVDD/1454 DVDD:13370 DVDD:13373 0.03348
rDVDD/1455 DVDD:13370 DVDD:13371 0.5625
rDVDD/1456 DVDD:13368 DVDD:15553 0.0292323
rDVDD/1457 DVDD:13367 DVDD:13370 0.03348
rDVDD/1458 DVDD:13367 DVDD:13368 0.5625
rDVDD/1459 DVDD:13365 DVDD:15548 0.0147047
rDVDD/1460 DVDD:13365 DVDD:13368 0.043937
rDVDD/1461 DVDD:13364 DVDD:13367 0.02232
rDVDD/1462 DVDD:13364 DVDD:13365 0.5625
rDVDD/1463 DVDD:13362 DVDD:15548 0.0512008
rDVDD/1464 DVDD:13361 DVDD:13364 0.03348
rDVDD/1465 DVDD:13361 DVDD:13362 0.5625
rDVDD/1466 DVDD:13359 DVDD:15543 0.0115157
rDVDD/1467 DVDD:13359 DVDD:13362 0.0659055
rDVDD/1468 DVDD:13358 DVDD:13361 0.03348
rDVDD/1469 DVDD:13358 DVDD:13359 0.5625
rDVDD/1470 DVDD:13356 DVDD:15539 0.0115157
rDVDD/1471 DVDD:13356 DVDD:15543 0.0324213
rDVDD/1472 DVDD:13355 DVDD:13358 0.02232
rDVDD/1473 DVDD:13355 DVDD:13356 0.5625
rDVDD/1474 DVDD:13348 DVDD:15533 0.028878
rDVDD/1475 DVDD:13347 DVDD:13348 0.75
rDVDD/1476 DVDD:13345 DVDD:13348 0.043937
rDVDD/1477 DVDD:13344 DVDD:13347 0.02232
rDVDD/1478 DVDD:13344 DVDD:13345 0.5625
rDVDD/1479 DVDD:13342 DVDD:13345 0.0659055
rDVDD/1480 DVDD:13341 DVDD:13344 0.03348
rDVDD/1481 DVDD:13341 DVDD:13342 0.5625
rDVDD/1482 DVDD:13339 DVDD:13342 0.043937
rDVDD/1483 DVDD:13338 DVDD:13341 0.02232
rDVDD/1484 DVDD:13338 DVDD:13339 0.5625
rDVDD/1485 DVDD:13336 DVDD:13339 0.0659055
rDVDD/1486 DVDD:13335 DVDD:13338 0.03348
rDVDD/1487 DVDD:13335 DVDD:13336 0.5625
rDVDD/1488 DVDD:13333 DVDD:13336 0.0659055
rDVDD/1489 DVDD:13332 DVDD:13335 0.03348
rDVDD/1490 DVDD:13332 DVDD:13333 0.5625
rDVDD/1491 DVDD:13330 DVDD:15523 0.0536811
rDVDD/1492 DVDD:13330 DVDD:13333 0.043937
rDVDD/1493 DVDD:13329 DVDD:13332 0.02232
rDVDD/1494 DVDD:13329 DVDD:13330 0.5625
rDVDD/1495 DVDD:13327 DVDD:15519 0.0536811
rDVDD/1496 DVDD:13327 DVDD:15523 0.0122244
rDVDD/1497 DVDD:13326 DVDD:13329 0.03348
rDVDD/1498 DVDD:13326 DVDD:13327 0.5625
rDVDD/1499 DVDD:13324 DVDD:15519 0.0122244
rDVDD/1500 DVDD:13323 DVDD:13326 0.03348
rDVDD/1501 DVDD:13323 DVDD:13324 0.5625
rDVDD/1502 DVDD:13321 DVDD:15514 0.0317126
rDVDD/1503 DVDD:13321 DVDD:13324 0.043937
rDVDD/1504 DVDD:13320 DVDD:13323 0.02232
rDVDD/1505 DVDD:13320 DVDD:13321 0.5625
rDVDD/1506 DVDD:13313 DVDD:15511 0.0965551
rDVDD/1507 DVDD:13313 DVDD:15436 0.3
rDVDD/1508 DVDD:13312 DVDD:13313 0.75
rDVDD/1509 DVDD:13310 DVDD:15504 0.0352559
rDVDD/1510 DVDD:13310 DVDD:13313 0.043937
rDVDD/1511 DVDD:13309 DVDD:13312 0.02232
rDVDD/1512 DVDD:13309 DVDD:13310 0.5625
rDVDD/1513 DVDD:13307 DVDD:15504 0.0306496
rDVDD/1514 DVDD:13306 DVDD:13309 0.03348
rDVDD/1515 DVDD:13306 DVDD:13307 0.5625
rDVDD/1516 DVDD:13304 DVDD:15499 0.0529724
rDVDD/1517 DVDD:13304 DVDD:13307 0.043937
rDVDD/1518 DVDD:13303 DVDD:13306 0.02232
rDVDD/1519 DVDD:13303 DVDD:13304 0.5625
rDVDD/1520 DVDD:13301 DVDD:15495 0.0310039
rDVDD/1521 DVDD:13301 DVDD:15499 0.0129331
rDVDD/1522 DVDD:13300 DVDD:13303 0.03348
rDVDD/1523 DVDD:13300 DVDD:13301 0.5625
rDVDD/1524 DVDD:13298 DVDD:15491 0.0310039
rDVDD/1525 DVDD:13298 DVDD:15495 0.0349016
rDVDD/1526 DVDD:13297 DVDD:13300 0.03348
rDVDD/1527 DVDD:13297 DVDD:13298 0.5625
rDVDD/1528 DVDD:13295 DVDD:15487 0.0749409
rDVDD/1529 DVDD:13295 DVDD:15491 0.0129331
rDVDD/1530 DVDD:13294 DVDD:13297 0.02232
rDVDD/1531 DVDD:13294 DVDD:13295 0.5625
rDVDD/1532 DVDD:13291 DVDD:13294 0.03348
rDVDD/1533 DVDD:13291 DVDD:15487 0.5625
rDVDD/1534 DVDD:13288 DVDD:13291 0.03348
rDVDD/1535 DVDD:13288 DVDD:15484 0.5625
rDVDD/1536 DVDD:13286 DVDD:15480 0.0529724
rDVDD/1537 DVDD:13286 DVDD:15484 0.0349016
rDVDD/1538 DVDD:13285 DVDD:13288 0.02232
rDVDD/1539 DVDD:13285 DVDD:13286 0.5625
rDVDD/1540 DVDD:13275 DVDD:13277 2.28827
rDVDD/1541 DVDD:13274 DVDD:13277 0.01944
rDVDD/1542 DVDD:13274 DVDD:13275 1.5
rDVDD/1543 DVDD:13272 DVDD:13275 0.0574016
rDVDD/1544 DVDD:13271 DVDD:13274 0.02916
rDVDD/1545 DVDD:13271 DVDD:13272 1.5
rDVDD/1546 DVDD:13269 DVDD:15211 0.0210827
rDVDD/1547 DVDD:13269 DVDD:13272 0.0574016
rDVDD/1548 DVDD:13268 DVDD:13271 0.02916
rDVDD/1549 DVDD:13268 DVDD:13269 1.5
rDVDD/1550 DVDD:13266 DVDD:15207 0.0295866
rDVDD/1551 DVDD:13266 DVDD:15211 0.0363189
rDVDD/1552 DVDD:13265 DVDD:13268 0.02916
rDVDD/1553 DVDD:13265 DVDD:13266 1.5
rDVDD/1554 DVDD:13263 DVDD:15207 0.027815
rDVDD/1555 DVDD:13262 DVDD:13265 0.02916
rDVDD/1556 DVDD:13262 DVDD:13263 1.5
rDVDD/1557 DVDD:13260 DVDD:15202 0.00265748
rDVDD/1558 DVDD:13260 DVDD:13263 0.0574016
rDVDD/1559 DVDD:13259 DVDD:13262 0.02916
rDVDD/1560 DVDD:13259 DVDD:13260 1.5
rDVDD/1561 DVDD:13257 DVDD:15202 0.0547441
rDVDD/1562 DVDD:13256 DVDD:13259 0.02916
rDVDD/1563 DVDD:13256 DVDD:13257 1.5
rDVDD/1564 DVDD:13254 DVDD:13257 0.0574016
rDVDD/1565 DVDD:13253 DVDD:13256 0.02916
rDVDD/1566 DVDD:13253 DVDD:13254 1.5
rDVDD/1567 DVDD:13251 DVDD:13254 0.0574016
rDVDD/1568 DVDD:13250 DVDD:13253 0.02916
rDVDD/1569 DVDD:13250 DVDD:13251 1.5
rDVDD/1570 DVDD:13243 DVDD:13251 0.201969
rDVDD/1571 DVDD:13242 DVDD:13243 2.25
rDVDD/1572 DVDD:13240 DVDD:13243 0.0382677
rDVDD/1573 DVDD:13239 DVDD:13242 0.01944
rDVDD/1574 DVDD:13239 DVDD:13240 1.5
rDVDD/1575 DVDD:13237 DVDD:13240 0.0574016
rDVDD/1576 DVDD:13236 DVDD:13239 0.02916
rDVDD/1577 DVDD:13236 DVDD:13237 1.5
rDVDD/1578 DVDD:13234 DVDD:13237 0.0574016
rDVDD/1579 DVDD:13233 DVDD:13236 0.02916
rDVDD/1580 DVDD:13233 DVDD:13234 1.5
rDVDD/1581 DVDD:13231 DVDD:13234 0.0574016
rDVDD/1582 DVDD:13230 DVDD:13233 0.02916
rDVDD/1583 DVDD:13230 DVDD:13231 1.5
rDVDD/1584 DVDD:13228 DVDD:13231 0.0574016
rDVDD/1585 DVDD:13227 DVDD:13230 0.02916
rDVDD/1586 DVDD:13227 DVDD:13228 1.5
rDVDD/1587 DVDD:13225 DVDD:13228 0.0574016
rDVDD/1588 DVDD:13224 DVDD:13227 0.02916
rDVDD/1589 DVDD:13224 DVDD:13225 1.5
rDVDD/1590 DVDD:13222 DVDD:13225 0.0574016
rDVDD/1591 DVDD:13221 DVDD:13224 0.02916
rDVDD/1592 DVDD:13221 DVDD:13222 1.5
rDVDD/1593 DVDD:13219 DVDD:13222 0.0574016
rDVDD/1594 DVDD:13218 DVDD:13221 0.02916
rDVDD/1595 DVDD:13218 DVDD:13219 1.5
rDVDD/1596 DVDD:13216 DVDD:13219 0.0574016
rDVDD/1597 DVDD:13215 DVDD:13218 0.02916
rDVDD/1598 DVDD:13215 DVDD:13216 1.5
rDVDD/1599 DVDD:13208 DVDD:13216 0.201969
rDVDD/1600 DVDD:13207 DVDD:13208 2.25
rDVDD/1601 DVDD:13205 DVDD:13208 0.0382677
rDVDD/1602 DVDD:13204 DVDD:13207 0.01944
rDVDD/1603 DVDD:13204 DVDD:13205 1.5
rDVDD/1604 DVDD:13202 DVDD:13205 0.0574016
rDVDD/1605 DVDD:13201 DVDD:13204 0.02916
rDVDD/1606 DVDD:13201 DVDD:13202 1.5
rDVDD/1607 DVDD:13199 DVDD:15182 0.0395079
rDVDD/1608 DVDD:13199 DVDD:13202 0.0574016
rDVDD/1609 DVDD:13198 DVDD:13201 0.02916
rDVDD/1610 DVDD:13198 DVDD:13199 1.5
rDVDD/1611 DVDD:13196 DVDD:15178 0.0480118
rDVDD/1612 DVDD:13196 DVDD:15182 0.0178937
rDVDD/1613 DVDD:13195 DVDD:13198 0.02916
rDVDD/1614 DVDD:13195 DVDD:13196 1.5
rDVDD/1615 DVDD:13193 DVDD:15178 0.00938976
rDVDD/1616 DVDD:13192 DVDD:13195 0.02916
rDVDD/1617 DVDD:13192 DVDD:13193 1.5
rDVDD/1618 DVDD:13190 DVDD:15173 0.0210827
rDVDD/1619 DVDD:13190 DVDD:13193 0.0574016
rDVDD/1620 DVDD:13189 DVDD:13192 0.02916
rDVDD/1621 DVDD:13189 DVDD:13190 1.5
rDVDD/1622 DVDD:13187 DVDD:15173 0.0363189
rDVDD/1623 DVDD:13186 DVDD:13189 0.02916
rDVDD/1624 DVDD:13186 DVDD:13187 1.5
rDVDD/1625 DVDD:13184 DVDD:13187 0.0574016
rDVDD/1626 DVDD:13183 DVDD:13186 0.02916
rDVDD/1627 DVDD:13183 DVDD:13184 1.5
rDVDD/1628 DVDD:13181 DVDD:13184 0.0574016
rDVDD/1629 DVDD:13180 DVDD:13183 0.02916
rDVDD/1630 DVDD:13180 DVDD:13181 1.5
rDVDD/1631 DVDD:13173 DVDD:15166 0.016122
rDVDD/1632 DVDD:13173 DVDD:13181 0.201969
rDVDD/1633 DVDD:13172 DVDD:13173 2.25
rDVDD/1634 DVDD:13170 DVDD:15162 0.0437598
rDVDD/1635 DVDD:13170 DVDD:15166 0.0221457
rDVDD/1636 DVDD:13169 DVDD:13172 0.01944
rDVDD/1637 DVDD:13169 DVDD:13170 1.5
rDVDD/1638 DVDD:13167 DVDD:15162 0.0136417
rDVDD/1639 DVDD:13166 DVDD:13169 0.02916
rDVDD/1640 DVDD:13166 DVDD:13167 1.5
rDVDD/1641 DVDD:13164 DVDD:15157 0.0168307
rDVDD/1642 DVDD:13164 DVDD:13167 0.0574016
rDVDD/1643 DVDD:13163 DVDD:13166 0.02916
rDVDD/1644 DVDD:13163 DVDD:13164 1.5
rDVDD/1645 DVDD:13161 DVDD:15157 0.0405709
rDVDD/1646 DVDD:13160 DVDD:13163 0.02916
rDVDD/1647 DVDD:13160 DVDD:13161 1.5
rDVDD/1648 DVDD:13158 DVDD:15152 0.0317126
rDVDD/1649 DVDD:13158 DVDD:13161 0.0574016
rDVDD/1650 DVDD:13157 DVDD:13160 0.02916
rDVDD/1651 DVDD:13157 DVDD:13158 1.5
rDVDD/1652 DVDD:13155 DVDD:15152 0.025689
rDVDD/1653 DVDD:13154 DVDD:13157 0.02916
rDVDD/1654 DVDD:13154 DVDD:13155 1.5
rDVDD/1655 DVDD:13152 DVDD:15147 0.00478346
rDVDD/1656 DVDD:13152 DVDD:13155 0.0574016
rDVDD/1657 DVDD:13151 DVDD:13154 0.02916
rDVDD/1658 DVDD:13151 DVDD:13152 1.5
rDVDD/1659 DVDD:13149 DVDD:15143 0.0132874
rDVDD/1660 DVDD:13149 DVDD:15147 0.0526181
rDVDD/1661 DVDD:13148 DVDD:13151 0.02916
rDVDD/1662 DVDD:13148 DVDD:13149 1.5
rDVDD/1663 DVDD:13146 DVDD:15139 0.0855709
rDVDD/1664 DVDD:13146 DVDD:15143 0.0441142
rDVDD/1665 DVDD:13145 DVDD:13148 0.02916
rDVDD/1666 DVDD:13145 DVDD:13146 1.5
rDVDD/1667 DVDD:13138 DVDD:15133 0.00655512
rDVDD/1668 DVDD:13137 DVDD:13138 2.25
rDVDD/1669 DVDD:13135 DVDD:15128 0.0430512
rDVDD/1670 DVDD:13135 DVDD:13138 0.0382677
rDVDD/1671 DVDD:13134 DVDD:13137 0.01944
rDVDD/1672 DVDD:13134 DVDD:13135 1.5
rDVDD/1673 DVDD:13132 DVDD:15128 0.0143504
rDVDD/1674 DVDD:13131 DVDD:13134 0.02916
rDVDD/1675 DVDD:13131 DVDD:13132 1.5
rDVDD/1676 DVDD:13129 DVDD:13132 0.0574016
rDVDD/1677 DVDD:13128 DVDD:13131 0.02916
rDVDD/1678 DVDD:13128 DVDD:13129 1.5
rDVDD/1679 DVDD:13126 DVDD:13129 0.0574016
rDVDD/1680 DVDD:13125 DVDD:13128 0.02916
rDVDD/1681 DVDD:13125 DVDD:13126 1.5
rDVDD/1682 DVDD:13123 DVDD:13126 0.0574016
rDVDD/1683 DVDD:13122 DVDD:13125 0.02916
rDVDD/1684 DVDD:13122 DVDD:13123 1.5
rDVDD/1685 DVDD:13120 DVDD:13123 0.0574016
rDVDD/1686 DVDD:13119 DVDD:13122 0.02916
rDVDD/1687 DVDD:13119 DVDD:13120 1.5
rDVDD/1688 DVDD:13117 DVDD:13120 0.0574016
rDVDD/1689 DVDD:13116 DVDD:13119 0.02916
rDVDD/1690 DVDD:13116 DVDD:13117 1.5
rDVDD/1691 DVDD:13114 DVDD:13117 0.0574016
rDVDD/1692 DVDD:13113 DVDD:13116 0.02916
rDVDD/1693 DVDD:13113 DVDD:13114 1.5
rDVDD/1694 DVDD:13111 DVDD:13114 0.0574016
rDVDD/1695 DVDD:13110 DVDD:13113 0.02916
rDVDD/1696 DVDD:13110 DVDD:13111 1.5
rDVDD/1697 DVDD:13103 DVDD:13111 0.201969
rDVDD/1698 DVDD:13102 DVDD:13103 2.25
rDVDD/1699 DVDD:13100 DVDD:13103 0.0382677
rDVDD/1700 DVDD:13099 DVDD:13102 0.01944
rDVDD/1701 DVDD:13099 DVDD:13100 1.5
rDVDD/1702 DVDD:13097 DVDD:13100 0.0574016
rDVDD/1703 DVDD:13096 DVDD:13099 0.02916
rDVDD/1704 DVDD:13096 DVDD:13097 1.5
rDVDD/1705 DVDD:13094 DVDD:13097 0.0574016
rDVDD/1706 DVDD:13093 DVDD:13096 0.02916
rDVDD/1707 DVDD:13093 DVDD:13094 1.5
rDVDD/1708 DVDD:13091 DVDD:13094 0.0574016
rDVDD/1709 DVDD:13090 DVDD:13093 0.02916
rDVDD/1710 DVDD:13090 DVDD:13091 1.5
rDVDD/1711 DVDD:13088 DVDD:13091 0.0574016
rDVDD/1712 DVDD:13087 DVDD:13090 0.02916
rDVDD/1713 DVDD:13087 DVDD:13088 1.5
rDVDD/1714 DVDD:13085 DVDD:13088 0.0574016
rDVDD/1715 DVDD:13084 DVDD:13087 0.02916
rDVDD/1716 DVDD:13084 DVDD:13085 1.5
rDVDD/1717 DVDD:13082 DVDD:13085 0.0574016
rDVDD/1718 DVDD:13081 DVDD:13084 0.02916
rDVDD/1719 DVDD:13081 DVDD:13082 1.5
rDVDD/1720 DVDD:13079 DVDD:13082 0.0574016
rDVDD/1721 DVDD:13078 DVDD:13081 0.02916
rDVDD/1722 DVDD:13078 DVDD:13079 1.5
rDVDD/1723 DVDD:13076 DVDD:15107 0.14687
rDVDD/1724 DVDD:13076 DVDD:13079 0.0574016
rDVDD/1725 DVDD:13075 DVDD:13078 0.02916
rDVDD/1726 DVDD:13075 DVDD:13076 1.5
rDVDD/1727 DVDD:13068 DVDD:15103 0.0108071
rDVDD/1728 DVDD:13068 DVDD:15107 0.0550984
rDVDD/1729 DVDD:13067 DVDD:13068 2.25
rDVDD/1730 DVDD:13065 DVDD:15103 0.0274606
rDVDD/1731 DVDD:13064 DVDD:13067 0.01944
rDVDD/1732 DVDD:13064 DVDD:13065 1.5
rDVDD/1733 DVDD:13062 DVDD:15098 0.00301181
rDVDD/1734 DVDD:13062 DVDD:13065 0.0574016
rDVDD/1735 DVDD:13061 DVDD:13064 0.02916
rDVDD/1736 DVDD:13061 DVDD:13062 1.5
rDVDD/1737 DVDD:13059 DVDD:15094 0.0115157
rDVDD/1738 DVDD:13059 DVDD:15098 0.0543898
rDVDD/1739 DVDD:13058 DVDD:13061 0.02916
rDVDD/1740 DVDD:13058 DVDD:13059 1.5
rDVDD/1741 DVDD:13056 DVDD:15090 0.0419882
rDVDD/1742 DVDD:13056 DVDD:15094 0.0458858
rDVDD/1743 DVDD:13055 DVDD:13058 0.02916
rDVDD/1744 DVDD:13055 DVDD:13056 1.5
rDVDD/1745 DVDD:13053 DVDD:15090 0.0154134
rDVDD/1746 DVDD:13052 DVDD:13055 0.02916
rDVDD/1747 DVDD:13052 DVDD:13053 1.5
rDVDD/1748 DVDD:13050 DVDD:15085 0.0150591
rDVDD/1749 DVDD:13050 DVDD:13053 0.0574016
rDVDD/1750 DVDD:13049 DVDD:13052 0.02916
rDVDD/1751 DVDD:13049 DVDD:13050 1.5
rDVDD/1752 DVDD:13047 DVDD:15085 0.0423425
rDVDD/1753 DVDD:13046 DVDD:13049 0.02916
rDVDD/1754 DVDD:13046 DVDD:13047 1.5
rDVDD/1755 DVDD:13044 DVDD:15080 0.028878
rDVDD/1756 DVDD:13044 DVDD:13047 0.0574016
rDVDD/1757 DVDD:13043 DVDD:13046 0.02916
rDVDD/1758 DVDD:13043 DVDD:13044 1.5
rDVDD/1759 DVDD:13041 DVDD:15076 0.0154134
rDVDD/1760 DVDD:13041 DVDD:15080 0.0285236
rDVDD/1761 DVDD:13040 DVDD:13043 0.02916
rDVDD/1762 DVDD:13040 DVDD:13041 1.5
rDVDD/1763 DVDD:13033 DVDD:15070 0.0327756
rDVDD/1764 DVDD:13032 DVDD:13033 2.25
rDVDD/1765 DVDD:13030 DVDD:13033 0.0382677
rDVDD/1766 DVDD:13029 DVDD:13032 0.01944
rDVDD/1767 DVDD:13029 DVDD:13030 1.5
rDVDD/1768 DVDD:13027 DVDD:13030 0.0574016
rDVDD/1769 DVDD:13026 DVDD:13029 0.02916
rDVDD/1770 DVDD:13026 DVDD:13027 1.5
rDVDD/1771 DVDD:13024 DVDD:13027 0.0574016
rDVDD/1772 DVDD:13023 DVDD:13026 0.02916
rDVDD/1773 DVDD:13023 DVDD:13024 1.5
rDVDD/1774 DVDD:13021 DVDD:13024 0.0574016
rDVDD/1775 DVDD:13020 DVDD:13023 0.02916
rDVDD/1776 DVDD:13020 DVDD:13021 1.5
rDVDD/1777 DVDD:13018 DVDD:13021 0.0574016
rDVDD/1778 DVDD:13017 DVDD:13020 0.02916
rDVDD/1779 DVDD:13017 DVDD:13018 1.5
rDVDD/1780 DVDD:13015 DVDD:15060 0.0540354
rDVDD/1781 DVDD:13015 DVDD:13018 0.0574016
rDVDD/1782 DVDD:13014 DVDD:13017 0.02916
rDVDD/1783 DVDD:13014 DVDD:13015 1.5
rDVDD/1784 DVDD:13012 DVDD:15060 0.00336614
rDVDD/1785 DVDD:13011 DVDD:13014 0.02916
rDVDD/1786 DVDD:13011 DVDD:13012 1.5
rDVDD/1787 DVDD:13009 DVDD:15055 0.0051378
rDVDD/1788 DVDD:13009 DVDD:13012 0.0574016
rDVDD/1789 DVDD:13008 DVDD:13011 0.02916
rDVDD/1790 DVDD:13008 DVDD:13009 1.5
rDVDD/1791 DVDD:13006 DVDD:15051 0.0356102
rDVDD/1792 DVDD:13006 DVDD:15055 0.0522638
rDVDD/1793 DVDD:13005 DVDD:13008 0.02916
rDVDD/1794 DVDD:13005 DVDD:13006 1.5
rDVDD/1795 DVDD:12998 DVDD:15045 0.0125787
rDVDD/1796 DVDD:12997 DVDD:12998 2.25
rDVDD/1797 DVDD:12995 DVDD:15040 0.0370276
rDVDD/1798 DVDD:12995 DVDD:12998 0.0382677
rDVDD/1799 DVDD:12994 DVDD:12997 0.01944
rDVDD/1800 DVDD:12994 DVDD:12995 1.5
rDVDD/1801 DVDD:12992 DVDD:15040 0.020374
rDVDD/1802 DVDD:12991 DVDD:12994 0.02916
rDVDD/1803 DVDD:12991 DVDD:12992 1.5
rDVDD/1804 DVDD:12989 DVDD:15035 0.0497835
rDVDD/1805 DVDD:12989 DVDD:12992 0.0574016
rDVDD/1806 DVDD:12988 DVDD:12991 0.02916
rDVDD/1807 DVDD:12988 DVDD:12989 1.5
rDVDD/1808 DVDD:12986 DVDD:15031 0.0363189
rDVDD/1809 DVDD:12986 DVDD:15035 0.00761811
rDVDD/1810 DVDD:12985 DVDD:12988 0.02916
rDVDD/1811 DVDD:12985 DVDD:12986 1.5
rDVDD/1812 DVDD:12983 DVDD:15027 0.0448228
rDVDD/1813 DVDD:12983 DVDD:15031 0.0210827
rDVDD/1814 DVDD:12982 DVDD:12985 0.02916
rDVDD/1815 DVDD:12982 DVDD:12983 1.5
rDVDD/1816 DVDD:12980 DVDD:15027 0.0125787
rDVDD/1817 DVDD:12979 DVDD:12982 0.02916
rDVDD/1818 DVDD:12979 DVDD:12980 1.5
rDVDD/1819 DVDD:12977 DVDD:15022 0.0178937
rDVDD/1820 DVDD:12977 DVDD:12980 0.0574016
rDVDD/1821 DVDD:12976 DVDD:12979 0.02916
rDVDD/1822 DVDD:12976 DVDD:12977 1.5
rDVDD/1823 DVDD:12974 DVDD:15018 0.0263976
rDVDD/1824 DVDD:12974 DVDD:15022 0.0395079
rDVDD/1825 DVDD:12973 DVDD:12976 0.02916
rDVDD/1826 DVDD:12973 DVDD:12974 1.5
rDVDD/1827 DVDD:12971 DVDD:15014 0.0568701
rDVDD/1828 DVDD:12971 DVDD:15018 0.0310039
rDVDD/1829 DVDD:12970 DVDD:12973 0.02916
rDVDD/1830 DVDD:12970 DVDD:12971 1.5
rDVDD/1831 DVDD:12960 DVDD:12962 2.28827
rDVDD/1832 DVDD:12959 DVDD:12962 0.01944
rDVDD/1833 DVDD:12959 DVDD:12960 1.5
rDVDD/1834 DVDD:12957 DVDD:12960 0.0574016
rDVDD/1835 DVDD:12956 DVDD:12959 0.02916
rDVDD/1836 DVDD:12956 DVDD:12957 1.5
rDVDD/1837 DVDD:12954 DVDD:14932 0.0210827
rDVDD/1838 DVDD:12954 DVDD:12957 0.0574016
rDVDD/1839 DVDD:12953 DVDD:12956 0.02916
rDVDD/1840 DVDD:12953 DVDD:12954 1.5
rDVDD/1841 DVDD:12951 DVDD:14928 0.0295866
rDVDD/1842 DVDD:12951 DVDD:14932 0.0363189
rDVDD/1843 DVDD:12950 DVDD:12953 0.02916
rDVDD/1844 DVDD:12950 DVDD:12951 1.5
rDVDD/1845 DVDD:12948 DVDD:14928 0.027815
rDVDD/1846 DVDD:12947 DVDD:12950 0.02916
rDVDD/1847 DVDD:12947 DVDD:12948 1.5
rDVDD/1848 DVDD:12945 DVDD:14923 0.00265748
rDVDD/1849 DVDD:12945 DVDD:12948 0.0574016
rDVDD/1850 DVDD:12944 DVDD:12947 0.02916
rDVDD/1851 DVDD:12944 DVDD:12945 1.5
rDVDD/1852 DVDD:12942 DVDD:14923 0.0547441
rDVDD/1853 DVDD:12941 DVDD:12944 0.02916
rDVDD/1854 DVDD:12941 DVDD:12942 1.5
rDVDD/1855 DVDD:12939 DVDD:12942 0.0574016
rDVDD/1856 DVDD:12938 DVDD:12941 0.02916
rDVDD/1857 DVDD:12938 DVDD:12939 1.5
rDVDD/1858 DVDD:12936 DVDD:12939 0.0574016
rDVDD/1859 DVDD:12935 DVDD:12938 0.02916
rDVDD/1860 DVDD:12935 DVDD:12936 1.5
rDVDD/1861 DVDD:12928 DVDD:12936 0.201969
rDVDD/1862 DVDD:12927 DVDD:12928 2.25
rDVDD/1863 DVDD:12925 DVDD:12928 0.0382677
rDVDD/1864 DVDD:12924 DVDD:12927 0.01944
rDVDD/1865 DVDD:12924 DVDD:12925 1.5
rDVDD/1866 DVDD:12922 DVDD:12925 0.0574016
rDVDD/1867 DVDD:12921 DVDD:12924 0.02916
rDVDD/1868 DVDD:12921 DVDD:12922 1.5
rDVDD/1869 DVDD:12919 DVDD:12922 0.0574016
rDVDD/1870 DVDD:12918 DVDD:12921 0.02916
rDVDD/1871 DVDD:12918 DVDD:12919 1.5
rDVDD/1872 DVDD:12916 DVDD:12919 0.0574016
rDVDD/1873 DVDD:12915 DVDD:12918 0.02916
rDVDD/1874 DVDD:12915 DVDD:12916 1.5
rDVDD/1875 DVDD:12913 DVDD:12916 0.0574016
rDVDD/1876 DVDD:12912 DVDD:12915 0.02916
rDVDD/1877 DVDD:12912 DVDD:12913 1.5
rDVDD/1878 DVDD:12910 DVDD:12913 0.0574016
rDVDD/1879 DVDD:12909 DVDD:12912 0.02916
rDVDD/1880 DVDD:12909 DVDD:12910 1.5
rDVDD/1881 DVDD:12907 DVDD:12910 0.0574016
rDVDD/1882 DVDD:12906 DVDD:12909 0.02916
rDVDD/1883 DVDD:12906 DVDD:12907 1.5
rDVDD/1884 DVDD:12904 DVDD:12907 0.0574016
rDVDD/1885 DVDD:12903 DVDD:12906 0.02916
rDVDD/1886 DVDD:12903 DVDD:12904 1.5
rDVDD/1887 DVDD:12901 DVDD:12904 0.0574016
rDVDD/1888 DVDD:12900 DVDD:12903 0.02916
rDVDD/1889 DVDD:12900 DVDD:12901 1.5
rDVDD/1890 DVDD:12893 DVDD:12901 0.201969
rDVDD/1891 DVDD:12892 DVDD:12893 2.25
rDVDD/1892 DVDD:12890 DVDD:12893 0.0382677
rDVDD/1893 DVDD:12889 DVDD:12892 0.01944
rDVDD/1894 DVDD:12889 DVDD:12890 1.5
rDVDD/1895 DVDD:12887 DVDD:12890 0.0574016
rDVDD/1896 DVDD:12886 DVDD:12889 0.02916
rDVDD/1897 DVDD:12886 DVDD:12887 1.5
rDVDD/1898 DVDD:12884 DVDD:14903 0.0395079
rDVDD/1899 DVDD:12884 DVDD:12887 0.0574016
rDVDD/1900 DVDD:12883 DVDD:12886 0.02916
rDVDD/1901 DVDD:12883 DVDD:12884 1.5
rDVDD/1902 DVDD:12881 DVDD:14899 0.0480118
rDVDD/1903 DVDD:12881 DVDD:14903 0.0178937
rDVDD/1904 DVDD:12880 DVDD:12883 0.02916
rDVDD/1905 DVDD:12880 DVDD:12881 1.5
rDVDD/1906 DVDD:12878 DVDD:14899 0.00938976
rDVDD/1907 DVDD:12877 DVDD:12880 0.02916
rDVDD/1908 DVDD:12877 DVDD:12878 1.5
rDVDD/1909 DVDD:12875 DVDD:14894 0.0210827
rDVDD/1910 DVDD:12875 DVDD:12878 0.0574016
rDVDD/1911 DVDD:12874 DVDD:12877 0.02916
rDVDD/1912 DVDD:12874 DVDD:12875 1.5
rDVDD/1913 DVDD:12872 DVDD:14894 0.0363189
rDVDD/1914 DVDD:12871 DVDD:12874 0.02916
rDVDD/1915 DVDD:12871 DVDD:12872 1.5
rDVDD/1916 DVDD:12869 DVDD:12872 0.0574016
rDVDD/1917 DVDD:12868 DVDD:12871 0.02916
rDVDD/1918 DVDD:12868 DVDD:12869 1.5
rDVDD/1919 DVDD:12866 DVDD:12869 0.0574016
rDVDD/1920 DVDD:12865 DVDD:12868 0.02916
rDVDD/1921 DVDD:12865 DVDD:12866 1.5
rDVDD/1922 DVDD:12858 DVDD:14887 0.016122
rDVDD/1923 DVDD:12858 DVDD:12866 0.201969
rDVDD/1924 DVDD:12857 DVDD:12858 2.25
rDVDD/1925 DVDD:12855 DVDD:14883 0.0217913
rDVDD/1926 DVDD:12855 DVDD:14887 0.0221457
rDVDD/1927 DVDD:12854 DVDD:12857 0.01944
rDVDD/1928 DVDD:12854 DVDD:12855 1.5
rDVDD/1929 DVDD:12852 DVDD:14879 0.0302953
rDVDD/1930 DVDD:12852 DVDD:14883 0.0356102
rDVDD/1931 DVDD:12851 DVDD:12854 0.02916
rDVDD/1932 DVDD:12851 DVDD:12852 1.5
rDVDD/1933 DVDD:12849 DVDD:14879 0.0271063
rDVDD/1934 DVDD:12848 DVDD:12851 0.02916
rDVDD/1935 DVDD:12848 DVDD:12849 1.5
rDVDD/1936 DVDD:12846 DVDD:14874 0.00336614
rDVDD/1937 DVDD:12846 DVDD:12849 0.0574016
rDVDD/1938 DVDD:12845 DVDD:12848 0.02916
rDVDD/1939 DVDD:12845 DVDD:12846 1.5
rDVDD/1940 DVDD:12843 DVDD:14870 0.0317126
rDVDD/1941 DVDD:12843 DVDD:14874 0.0540354
rDVDD/1942 DVDD:12842 DVDD:12845 0.02916
rDVDD/1943 DVDD:12842 DVDD:12843 1.5
rDVDD/1944 DVDD:12840 DVDD:14870 0.025689
rDVDD/1945 DVDD:12839 DVDD:12842 0.02916
rDVDD/1946 DVDD:12839 DVDD:12840 1.5
rDVDD/1947 DVDD:12837 DVDD:14865 0.00478346
rDVDD/1948 DVDD:12837 DVDD:12840 0.0574016
rDVDD/1949 DVDD:12836 DVDD:12839 0.02916
rDVDD/1950 DVDD:12836 DVDD:12837 1.5
rDVDD/1951 DVDD:12834 DVDD:14861 0.0132874
rDVDD/1952 DVDD:12834 DVDD:14865 0.0526181
rDVDD/1953 DVDD:12833 DVDD:12836 0.02916
rDVDD/1954 DVDD:12833 DVDD:12834 1.5
rDVDD/1955 DVDD:12831 DVDD:14857 0.0855709
rDVDD/1956 DVDD:12831 DVDD:14861 0.0441142
rDVDD/1957 DVDD:12830 DVDD:12833 0.02916
rDVDD/1958 DVDD:12830 DVDD:12831 1.5
rDVDD/1959 DVDD:12823 DVDD:14850 0.0154134
rDVDD/1960 DVDD:12823 DVDD:14854 0.0504921
rDVDD/1961 DVDD:12822 DVDD:12823 2.25
rDVDD/1962 DVDD:12820 DVDD:14846 0.0430512
rDVDD/1963 DVDD:12820 DVDD:14850 0.0228543
rDVDD/1964 DVDD:12819 DVDD:12822 0.01944
rDVDD/1965 DVDD:12819 DVDD:12820 1.5
rDVDD/1966 DVDD:12817 DVDD:14846 0.0143504
rDVDD/1967 DVDD:12816 DVDD:12819 0.02916
rDVDD/1968 DVDD:12816 DVDD:12817 1.5
rDVDD/1969 DVDD:12814 DVDD:12817 0.0574016
rDVDD/1970 DVDD:12813 DVDD:12816 0.02916
rDVDD/1971 DVDD:12813 DVDD:12814 1.5
rDVDD/1972 DVDD:12811 DVDD:12814 0.0574016
rDVDD/1973 DVDD:12810 DVDD:12813 0.02916
rDVDD/1974 DVDD:12810 DVDD:12811 1.5
rDVDD/1975 DVDD:12808 DVDD:12811 0.0574016
rDVDD/1976 DVDD:12807 DVDD:12810 0.02916
rDVDD/1977 DVDD:12807 DVDD:12808 1.5
rDVDD/1978 DVDD:12805 DVDD:12808 0.0574016
rDVDD/1979 DVDD:12804 DVDD:12807 0.02916
rDVDD/1980 DVDD:12804 DVDD:12805 1.5
rDVDD/1981 DVDD:12802 DVDD:12805 0.0574016
rDVDD/1982 DVDD:12801 DVDD:12804 0.02916
rDVDD/1983 DVDD:12801 DVDD:12802 1.5
rDVDD/1984 DVDD:12799 DVDD:12802 0.0574016
rDVDD/1985 DVDD:12798 DVDD:12801 0.02916
rDVDD/1986 DVDD:12798 DVDD:12799 1.5
rDVDD/1987 DVDD:12796 DVDD:12799 0.0574016
rDVDD/1988 DVDD:12795 DVDD:12798 0.02916
rDVDD/1989 DVDD:12795 DVDD:12796 1.5
rDVDD/1990 DVDD:12788 DVDD:12796 0.201969
rDVDD/1991 DVDD:12787 DVDD:12788 2.25
rDVDD/1992 DVDD:12785 DVDD:12788 0.0382677
rDVDD/1993 DVDD:12784 DVDD:12787 0.01944
rDVDD/1994 DVDD:12784 DVDD:12785 1.5
rDVDD/1995 DVDD:12782 DVDD:12785 0.0574016
rDVDD/1996 DVDD:12781 DVDD:12784 0.02916
rDVDD/1997 DVDD:12781 DVDD:12782 1.5
rDVDD/1998 DVDD:12779 DVDD:12782 0.0574016
rDVDD/1999 DVDD:12778 DVDD:12781 0.02916
rDVDD/2000 DVDD:12778 DVDD:12779 1.5
rDVDD/2001 DVDD:12776 DVDD:12779 0.0574016
rDVDD/2002 DVDD:12775 DVDD:12778 0.02916
rDVDD/2003 DVDD:12775 DVDD:12776 1.5
rDVDD/2004 DVDD:12773 DVDD:12776 0.0574016
rDVDD/2005 DVDD:12772 DVDD:12775 0.02916
rDVDD/2006 DVDD:12772 DVDD:12773 1.5
rDVDD/2007 DVDD:12770 DVDD:12773 0.0574016
rDVDD/2008 DVDD:12769 DVDD:12772 0.02916
rDVDD/2009 DVDD:12769 DVDD:12770 1.5
rDVDD/2010 DVDD:12767 DVDD:12770 0.0574016
rDVDD/2011 DVDD:12766 DVDD:12769 0.02916
rDVDD/2012 DVDD:12766 DVDD:12767 1.5
rDVDD/2013 DVDD:12764 DVDD:12767 0.0574016
rDVDD/2014 DVDD:12763 DVDD:12766 0.02916
rDVDD/2015 DVDD:12763 DVDD:12764 1.5
rDVDD/2016 DVDD:12761 DVDD:14825 0.14687
rDVDD/2017 DVDD:12761 DVDD:12764 0.0574016
rDVDD/2018 DVDD:12760 DVDD:12763 0.02916
rDVDD/2019 DVDD:12760 DVDD:12761 1.5
rDVDD/2020 DVDD:12753 DVDD:14821 0.0108071
rDVDD/2021 DVDD:12753 DVDD:14825 0.0550984
rDVDD/2022 DVDD:12752 DVDD:12753 2.25
rDVDD/2023 DVDD:12750 DVDD:14821 0.0274606
rDVDD/2024 DVDD:12749 DVDD:12752 0.01944
rDVDD/2025 DVDD:12749 DVDD:12750 1.5
rDVDD/2026 DVDD:12747 DVDD:14816 0.00301181
rDVDD/2027 DVDD:12747 DVDD:12750 0.0574016
rDVDD/2028 DVDD:12746 DVDD:12749 0.02916
rDVDD/2029 DVDD:12746 DVDD:12747 1.5
rDVDD/2030 DVDD:12744 DVDD:14812 0.0115157
rDVDD/2031 DVDD:12744 DVDD:14816 0.0543898
rDVDD/2032 DVDD:12743 DVDD:12746 0.02916
rDVDD/2033 DVDD:12743 DVDD:12744 1.5
rDVDD/2034 DVDD:12741 DVDD:14808 0.0419882
rDVDD/2035 DVDD:12741 DVDD:14812 0.0458858
rDVDD/2036 DVDD:12740 DVDD:12743 0.02916
rDVDD/2037 DVDD:12740 DVDD:12741 1.5
rDVDD/2038 DVDD:12738 DVDD:14804 0.0504921
rDVDD/2039 DVDD:12738 DVDD:14808 0.0154134
rDVDD/2040 DVDD:12737 DVDD:12740 0.02916
rDVDD/2041 DVDD:12737 DVDD:12738 1.5
rDVDD/2042 DVDD:12735 DVDD:14804 0.00690945
rDVDD/2043 DVDD:12734 DVDD:12737 0.02916
rDVDD/2044 DVDD:12734 DVDD:12735 1.5
rDVDD/2045 DVDD:12732 DVDD:14799 0.023563
rDVDD/2046 DVDD:12732 DVDD:12735 0.0574016
rDVDD/2047 DVDD:12731 DVDD:12734 0.02916
rDVDD/2048 DVDD:12731 DVDD:12732 1.5
rDVDD/2049 DVDD:12729 DVDD:14799 0.0338386
rDVDD/2050 DVDD:12728 DVDD:12731 0.02916
rDVDD/2051 DVDD:12728 DVDD:12729 1.5
rDVDD/2052 DVDD:12726 DVDD:14794 0.0154134
rDVDD/2053 DVDD:12726 DVDD:12729 0.0574016
rDVDD/2054 DVDD:12725 DVDD:12728 0.02916
rDVDD/2055 DVDD:12725 DVDD:12726 1.5
rDVDD/2056 DVDD:12718 DVDD:14788 0.0327756
rDVDD/2057 DVDD:12717 DVDD:12718 2.25
rDVDD/2058 DVDD:12715 DVDD:12718 0.0382677
rDVDD/2059 DVDD:12714 DVDD:12717 0.01944
rDVDD/2060 DVDD:12714 DVDD:12715 1.5
rDVDD/2061 DVDD:12712 DVDD:12715 0.0574016
rDVDD/2062 DVDD:12711 DVDD:12714 0.02916
rDVDD/2063 DVDD:12711 DVDD:12712 1.5
rDVDD/2064 DVDD:12709 DVDD:12712 0.0574016
rDVDD/2065 DVDD:12708 DVDD:12711 0.02916
rDVDD/2066 DVDD:12708 DVDD:12709 1.5
rDVDD/2067 DVDD:12706 DVDD:12709 0.0574016
rDVDD/2068 DVDD:12705 DVDD:12708 0.02916
rDVDD/2069 DVDD:12705 DVDD:12706 1.5
rDVDD/2070 DVDD:12703 DVDD:12706 0.0574016
rDVDD/2071 DVDD:12702 DVDD:12705 0.02916
rDVDD/2072 DVDD:12702 DVDD:12703 1.5
rDVDD/2073 DVDD:12700 DVDD:14778 0.0100984
rDVDD/2074 DVDD:12700 DVDD:12703 0.0574016
rDVDD/2075 DVDD:12699 DVDD:12702 0.02916
rDVDD/2076 DVDD:12699 DVDD:12700 1.5
rDVDD/2077 DVDD:12697 DVDD:14774 0.0186024
rDVDD/2078 DVDD:12697 DVDD:14778 0.0473032
rDVDD/2079 DVDD:12696 DVDD:12699 0.02916
rDVDD/2080 DVDD:12696 DVDD:12697 1.5
rDVDD/2081 DVDD:12694 DVDD:14770 0.0490748
rDVDD/2082 DVDD:12694 DVDD:14774 0.0387992
rDVDD/2083 DVDD:12693 DVDD:12696 0.02916
rDVDD/2084 DVDD:12693 DVDD:12694 1.5
rDVDD/2085 DVDD:12691 DVDD:14766 0.0575787
rDVDD/2086 DVDD:12691 DVDD:14770 0.00832677
rDVDD/2087 DVDD:12690 DVDD:12693 0.02916
rDVDD/2088 DVDD:12690 DVDD:12691 1.5
rDVDD/2089 DVDD:12683 DVDD:14759 0.00938976
rDVDD/2090 DVDD:12683 DVDD:14763 0.0565157
rDVDD/2091 DVDD:12682 DVDD:12683 2.25
rDVDD/2092 DVDD:12680 DVDD:14759 0.028878
rDVDD/2093 DVDD:12679 DVDD:12682 0.01944
rDVDD/2094 DVDD:12679 DVDD:12680 1.5
rDVDD/2095 DVDD:12677 DVDD:14754 0.00159449
rDVDD/2096 DVDD:12677 DVDD:12680 0.0574016
rDVDD/2097 DVDD:12676 DVDD:12679 0.02916
rDVDD/2098 DVDD:12676 DVDD:12677 1.5
rDVDD/2099 DVDD:12674 DVDD:14750 0.0497835
rDVDD/2100 DVDD:12674 DVDD:14754 0.0558071
rDVDD/2101 DVDD:12673 DVDD:12676 0.02916
rDVDD/2102 DVDD:12673 DVDD:12674 1.5
rDVDD/2103 DVDD:12671 DVDD:14750 0.00761811
rDVDD/2104 DVDD:12670 DVDD:12673 0.02916
rDVDD/2105 DVDD:12670 DVDD:12671 1.5
rDVDD/2106 DVDD:12668 DVDD:14745 0.0228543
rDVDD/2107 DVDD:12668 DVDD:12671 0.0574016
rDVDD/2108 DVDD:12667 DVDD:12670 0.02916
rDVDD/2109 DVDD:12667 DVDD:12668 1.5
rDVDD/2110 DVDD:12665 DVDD:14741 0.0313583
rDVDD/2111 DVDD:12665 DVDD:14745 0.0345472
rDVDD/2112 DVDD:12664 DVDD:12667 0.02916
rDVDD/2113 DVDD:12664 DVDD:12665 1.5
rDVDD/2114 DVDD:12662 DVDD:14741 0.0260433
rDVDD/2115 DVDD:12661 DVDD:12664 0.02916
rDVDD/2116 DVDD:12661 DVDD:12662 1.5
rDVDD/2117 DVDD:12659 DVDD:14736 0.00442913
rDVDD/2118 DVDD:12659 DVDD:12662 0.0574016
rDVDD/2119 DVDD:12658 DVDD:12661 0.02916
rDVDD/2120 DVDD:12658 DVDD:12659 1.5
rDVDD/2121 DVDD:12656 DVDD:14732 0.0129331
rDVDD/2122 DVDD:12656 DVDD:14736 0.0529724
rDVDD/2123 DVDD:12655 DVDD:12658 0.02916
rDVDD/2124 DVDD:12655 DVDD:12656 1.5
rDVDD/2125 DVDD:12645 DVDD:12647 2.28827
rDVDD/2126 DVDD:12644 DVDD:12647 0.01944
rDVDD/2127 DVDD:12644 DVDD:12645 1.5
rDVDD/2128 DVDD:12642 DVDD:12645 0.0574016
rDVDD/2129 DVDD:12641 DVDD:12644 0.02916
rDVDD/2130 DVDD:12641 DVDD:12642 1.5
rDVDD/2131 DVDD:12639 DVDD:14647 0.0210827
rDVDD/2132 DVDD:12639 DVDD:12642 0.0574016
rDVDD/2133 DVDD:12638 DVDD:12641 0.02916
rDVDD/2134 DVDD:12638 DVDD:12639 1.5
rDVDD/2135 DVDD:12636 DVDD:14643 0.0295866
rDVDD/2136 DVDD:12636 DVDD:14647 0.0363189
rDVDD/2137 DVDD:12635 DVDD:12638 0.02916
rDVDD/2138 DVDD:12635 DVDD:12636 1.5
rDVDD/2139 DVDD:12633 DVDD:14643 0.027815
rDVDD/2140 DVDD:12632 DVDD:12635 0.02916
rDVDD/2141 DVDD:12632 DVDD:12633 1.5
rDVDD/2142 DVDD:12630 DVDD:14638 0.00265748
rDVDD/2143 DVDD:12630 DVDD:12633 0.0574016
rDVDD/2144 DVDD:12629 DVDD:12632 0.02916
rDVDD/2145 DVDD:12629 DVDD:12630 1.5
rDVDD/2146 DVDD:12627 DVDD:14638 0.0547441
rDVDD/2147 DVDD:12626 DVDD:12629 0.02916
rDVDD/2148 DVDD:12626 DVDD:12627 1.5
rDVDD/2149 DVDD:12624 DVDD:12627 0.0574016
rDVDD/2150 DVDD:12623 DVDD:12626 0.02916
rDVDD/2151 DVDD:12623 DVDD:12624 1.5
rDVDD/2152 DVDD:12621 DVDD:12624 0.0574016
rDVDD/2153 DVDD:12620 DVDD:12623 0.02916
rDVDD/2154 DVDD:12620 DVDD:12621 1.5
rDVDD/2155 DVDD:12613 DVDD:12621 0.201969
rDVDD/2156 DVDD:12612 DVDD:12613 2.25
rDVDD/2157 DVDD:12610 DVDD:12613 0.0382677
rDVDD/2158 DVDD:12609 DVDD:12612 0.01944
rDVDD/2159 DVDD:12609 DVDD:12610 1.5
rDVDD/2160 DVDD:12607 DVDD:12610 0.0574016
rDVDD/2161 DVDD:12606 DVDD:12609 0.02916
rDVDD/2162 DVDD:12606 DVDD:12607 1.5
rDVDD/2163 DVDD:12604 DVDD:12607 0.0574016
rDVDD/2164 DVDD:12603 DVDD:12606 0.02916
rDVDD/2165 DVDD:12603 DVDD:12604 1.5
rDVDD/2166 DVDD:12601 DVDD:12604 0.0574016
rDVDD/2167 DVDD:12600 DVDD:12603 0.02916
rDVDD/2168 DVDD:12600 DVDD:12601 1.5
rDVDD/2169 DVDD:12598 DVDD:12601 0.0574016
rDVDD/2170 DVDD:12597 DVDD:12600 0.02916
rDVDD/2171 DVDD:12597 DVDD:12598 1.5
rDVDD/2172 DVDD:12595 DVDD:12598 0.0574016
rDVDD/2173 DVDD:12594 DVDD:12597 0.02916
rDVDD/2174 DVDD:12594 DVDD:12595 1.5
rDVDD/2175 DVDD:12592 DVDD:12595 0.0574016
rDVDD/2176 DVDD:12591 DVDD:12594 0.02916
rDVDD/2177 DVDD:12591 DVDD:12592 1.5
rDVDD/2178 DVDD:12589 DVDD:12592 0.0574016
rDVDD/2179 DVDD:12588 DVDD:12591 0.02916
rDVDD/2180 DVDD:12588 DVDD:12589 1.5
rDVDD/2181 DVDD:12586 DVDD:12589 0.0574016
rDVDD/2182 DVDD:12585 DVDD:12588 0.02916
rDVDD/2183 DVDD:12585 DVDD:12586 1.5
rDVDD/2184 DVDD:12578 DVDD:12586 0.201969
rDVDD/2185 DVDD:12577 DVDD:12578 2.25
rDVDD/2186 DVDD:12575 DVDD:12578 0.0382677
rDVDD/2187 DVDD:12574 DVDD:12577 0.01944
rDVDD/2188 DVDD:12574 DVDD:12575 1.5
rDVDD/2189 DVDD:12572 DVDD:12575 0.0574016
rDVDD/2190 DVDD:12571 DVDD:12574 0.02916
rDVDD/2191 DVDD:12571 DVDD:12572 1.5
rDVDD/2192 DVDD:12569 DVDD:14618 0.0395079
rDVDD/2193 DVDD:12569 DVDD:12572 0.0574016
rDVDD/2194 DVDD:12568 DVDD:12571 0.02916
rDVDD/2195 DVDD:12568 DVDD:12569 1.5
rDVDD/2196 DVDD:12566 DVDD:14614 0.0480118
rDVDD/2197 DVDD:12566 DVDD:14618 0.0178937
rDVDD/2198 DVDD:12565 DVDD:12568 0.02916
rDVDD/2199 DVDD:12565 DVDD:12566 1.5
rDVDD/2200 DVDD:12563 DVDD:14614 0.00938976
rDVDD/2201 DVDD:12562 DVDD:12565 0.02916
rDVDD/2202 DVDD:12562 DVDD:12563 1.5
rDVDD/2203 DVDD:12560 DVDD:14609 0.0210827
rDVDD/2204 DVDD:12560 DVDD:12563 0.0574016
rDVDD/2205 DVDD:12559 DVDD:12562 0.02916
rDVDD/2206 DVDD:12559 DVDD:12560 1.5
rDVDD/2207 DVDD:12557 DVDD:14609 0.0363189
rDVDD/2208 DVDD:12556 DVDD:12559 0.02916
rDVDD/2209 DVDD:12556 DVDD:12557 1.5
rDVDD/2210 DVDD:12554 DVDD:12557 0.0574016
rDVDD/2211 DVDD:12553 DVDD:12556 0.02916
rDVDD/2212 DVDD:12553 DVDD:12554 1.5
rDVDD/2213 DVDD:12551 DVDD:12554 0.0574016
rDVDD/2214 DVDD:12550 DVDD:12553 0.02916
rDVDD/2215 DVDD:12550 DVDD:12551 1.5
rDVDD/2216 DVDD:12543 DVDD:14602 0.016122
rDVDD/2217 DVDD:12543 DVDD:12551 0.201969
rDVDD/2218 DVDD:12542 DVDD:12543 2.25
rDVDD/2219 DVDD:12540 DVDD:14598 0.0217913
rDVDD/2220 DVDD:12540 DVDD:14602 0.0221457
rDVDD/2221 DVDD:12539 DVDD:12542 0.01944
rDVDD/2222 DVDD:12539 DVDD:12540 1.5
rDVDD/2223 DVDD:12537 DVDD:14594 0.0302953
rDVDD/2224 DVDD:12537 DVDD:14598 0.0356102
rDVDD/2225 DVDD:12536 DVDD:12539 0.02916
rDVDD/2226 DVDD:12536 DVDD:12537 1.5
rDVDD/2227 DVDD:12534 DVDD:14594 0.0271063
rDVDD/2228 DVDD:12533 DVDD:12536 0.02916
rDVDD/2229 DVDD:12533 DVDD:12534 1.5
rDVDD/2230 DVDD:12531 DVDD:14589 0.00336614
rDVDD/2231 DVDD:12531 DVDD:12534 0.0574016
rDVDD/2232 DVDD:12530 DVDD:12533 0.02916
rDVDD/2233 DVDD:12530 DVDD:12531 1.5
rDVDD/2234 DVDD:12528 DVDD:14585 0.0317126
rDVDD/2235 DVDD:12528 DVDD:14589 0.0540354
rDVDD/2236 DVDD:12527 DVDD:12530 0.02916
rDVDD/2237 DVDD:12527 DVDD:12528 1.5
rDVDD/2238 DVDD:12525 DVDD:14585 0.025689
rDVDD/2239 DVDD:12524 DVDD:12527 0.02916
rDVDD/2240 DVDD:12524 DVDD:12525 1.5
rDVDD/2241 DVDD:12522 DVDD:14580 0.00478346
rDVDD/2242 DVDD:12522 DVDD:12525 0.0574016
rDVDD/2243 DVDD:12521 DVDD:12524 0.02916
rDVDD/2244 DVDD:12521 DVDD:12522 1.5
rDVDD/2245 DVDD:12519 DVDD:14576 0.0132874
rDVDD/2246 DVDD:12519 DVDD:14580 0.0526181
rDVDD/2247 DVDD:12518 DVDD:12521 0.02916
rDVDD/2248 DVDD:12518 DVDD:12519 1.5
rDVDD/2249 DVDD:12516 DVDD:14572 0.0855709
rDVDD/2250 DVDD:12516 DVDD:14576 0.0441142
rDVDD/2251 DVDD:12515 DVDD:12518 0.02916
rDVDD/2252 DVDD:12515 DVDD:12516 1.5
rDVDD/2253 DVDD:12508 DVDD:14565 0.0154134
rDVDD/2254 DVDD:12508 DVDD:14569 0.0504921
rDVDD/2255 DVDD:12507 DVDD:12508 2.25
rDVDD/2256 DVDD:12505 DVDD:14561 0.0430512
rDVDD/2257 DVDD:12505 DVDD:14565 0.0228543
rDVDD/2258 DVDD:12504 DVDD:12507 0.01944
rDVDD/2259 DVDD:12504 DVDD:12505 1.5
rDVDD/2260 DVDD:12502 DVDD:14561 0.0143504
rDVDD/2261 DVDD:12501 DVDD:12504 0.02916
rDVDD/2262 DVDD:12501 DVDD:12502 1.5
rDVDD/2263 DVDD:12499 DVDD:12502 0.0574016
rDVDD/2264 DVDD:12498 DVDD:12501 0.02916
rDVDD/2265 DVDD:12498 DVDD:12499 1.5
rDVDD/2266 DVDD:12496 DVDD:12499 0.0574016
rDVDD/2267 DVDD:12495 DVDD:12498 0.02916
rDVDD/2268 DVDD:12495 DVDD:12496 1.5
rDVDD/2269 DVDD:12493 DVDD:12496 0.0574016
rDVDD/2270 DVDD:12492 DVDD:12495 0.02916
rDVDD/2271 DVDD:12492 DVDD:12493 1.5
rDVDD/2272 DVDD:12490 DVDD:12493 0.0574016
rDVDD/2273 DVDD:12489 DVDD:12492 0.02916
rDVDD/2274 DVDD:12489 DVDD:12490 1.5
rDVDD/2275 DVDD:12487 DVDD:12490 0.0574016
rDVDD/2276 DVDD:12486 DVDD:12489 0.02916
rDVDD/2277 DVDD:12486 DVDD:12487 1.5
rDVDD/2278 DVDD:12484 DVDD:12487 0.0574016
rDVDD/2279 DVDD:12483 DVDD:12486 0.02916
rDVDD/2280 DVDD:12483 DVDD:12484 1.5
rDVDD/2281 DVDD:12481 DVDD:12484 0.0574016
rDVDD/2282 DVDD:12480 DVDD:12483 0.02916
rDVDD/2283 DVDD:12480 DVDD:12481 1.5
rDVDD/2284 DVDD:12473 DVDD:12481 0.201969
rDVDD/2285 DVDD:12472 DVDD:12473 2.25
rDVDD/2286 DVDD:12470 DVDD:12473 0.0382677
rDVDD/2287 DVDD:12469 DVDD:12472 0.01944
rDVDD/2288 DVDD:12469 DVDD:12470 1.5
rDVDD/2289 DVDD:12467 DVDD:12470 0.0574016
rDVDD/2290 DVDD:12466 DVDD:12469 0.02916
rDVDD/2291 DVDD:12466 DVDD:12467 1.5
rDVDD/2292 DVDD:12464 DVDD:12467 0.0574016
rDVDD/2293 DVDD:12463 DVDD:12466 0.02916
rDVDD/2294 DVDD:12463 DVDD:12464 1.5
rDVDD/2295 DVDD:12461 DVDD:12464 0.0574016
rDVDD/2296 DVDD:12460 DVDD:12463 0.02916
rDVDD/2297 DVDD:12460 DVDD:12461 1.5
rDVDD/2298 DVDD:12458 DVDD:12461 0.0574016
rDVDD/2299 DVDD:12457 DVDD:12460 0.02916
rDVDD/2300 DVDD:12457 DVDD:12458 1.5
rDVDD/2301 DVDD:12455 DVDD:12458 0.0574016
rDVDD/2302 DVDD:12454 DVDD:12457 0.02916
rDVDD/2303 DVDD:12454 DVDD:12455 1.5
rDVDD/2304 DVDD:12452 DVDD:12455 0.0574016
rDVDD/2305 DVDD:12451 DVDD:12454 0.02916
rDVDD/2306 DVDD:12451 DVDD:12452 1.5
rDVDD/2307 DVDD:12449 DVDD:12452 0.0574016
rDVDD/2308 DVDD:12448 DVDD:12451 0.02916
rDVDD/2309 DVDD:12448 DVDD:12449 1.5
rDVDD/2310 DVDD:12446 DVDD:14540 0.14687
rDVDD/2311 DVDD:12446 DVDD:12449 0.0574016
rDVDD/2312 DVDD:12445 DVDD:12448 0.02916
rDVDD/2313 DVDD:12445 DVDD:12446 1.5
rDVDD/2314 DVDD:12438 DVDD:14536 0.0108071
rDVDD/2315 DVDD:12438 DVDD:14540 0.0550984
rDVDD/2316 DVDD:12437 DVDD:12438 2.25
rDVDD/2317 DVDD:12435 DVDD:14536 0.0274606
rDVDD/2318 DVDD:12434 DVDD:12437 0.01944
rDVDD/2319 DVDD:12434 DVDD:12435 1.5
rDVDD/2320 DVDD:12432 DVDD:14531 0.00301181
rDVDD/2321 DVDD:12432 DVDD:12435 0.0574016
rDVDD/2322 DVDD:12431 DVDD:12434 0.02916
rDVDD/2323 DVDD:12431 DVDD:12432 1.5
rDVDD/2324 DVDD:12429 DVDD:14527 0.0115157
rDVDD/2325 DVDD:12429 DVDD:14531 0.0543898
rDVDD/2326 DVDD:12428 DVDD:12431 0.02916
rDVDD/2327 DVDD:12428 DVDD:12429 1.5
rDVDD/2328 DVDD:12426 DVDD:14523 0.0419882
rDVDD/2329 DVDD:12426 DVDD:14527 0.0458858
rDVDD/2330 DVDD:12425 DVDD:12428 0.02916
rDVDD/2331 DVDD:12425 DVDD:12426 1.5
rDVDD/2332 DVDD:12423 DVDD:14519 0.0504921
rDVDD/2333 DVDD:12423 DVDD:14523 0.0154134
rDVDD/2334 DVDD:12422 DVDD:12425 0.02916
rDVDD/2335 DVDD:12422 DVDD:12423 1.5
rDVDD/2336 DVDD:12420 DVDD:14519 0.00690945
rDVDD/2337 DVDD:12419 DVDD:12422 0.02916
rDVDD/2338 DVDD:12419 DVDD:12420 1.5
rDVDD/2339 DVDD:12417 DVDD:14514 0.023563
rDVDD/2340 DVDD:12417 DVDD:12420 0.0574016
rDVDD/2341 DVDD:12416 DVDD:12419 0.02916
rDVDD/2342 DVDD:12416 DVDD:12417 1.5
rDVDD/2343 DVDD:12414 DVDD:14514 0.0338386
rDVDD/2344 DVDD:12413 DVDD:12416 0.02916
rDVDD/2345 DVDD:12413 DVDD:12414 1.5
rDVDD/2346 DVDD:12411 DVDD:14509 0.0154134
rDVDD/2347 DVDD:12411 DVDD:12414 0.0574016
rDVDD/2348 DVDD:12410 DVDD:12413 0.02916
rDVDD/2349 DVDD:12410 DVDD:12411 1.5
rDVDD/2350 DVDD:12403 DVDD:14503 0.0327756
rDVDD/2351 DVDD:12402 DVDD:12403 2.25
rDVDD/2352 DVDD:12400 DVDD:12403 0.0382677
rDVDD/2353 DVDD:12399 DVDD:12402 0.01944
rDVDD/2354 DVDD:12399 DVDD:12400 1.5
rDVDD/2355 DVDD:12397 DVDD:12400 0.0574016
rDVDD/2356 DVDD:12396 DVDD:12399 0.02916
rDVDD/2357 DVDD:12396 DVDD:12397 1.5
rDVDD/2358 DVDD:12394 DVDD:12397 0.0574016
rDVDD/2359 DVDD:12393 DVDD:12396 0.02916
rDVDD/2360 DVDD:12393 DVDD:12394 1.5
rDVDD/2361 DVDD:12391 DVDD:12394 0.0574016
rDVDD/2362 DVDD:12390 DVDD:12393 0.02916
rDVDD/2363 DVDD:12390 DVDD:12391 1.5
rDVDD/2364 DVDD:12388 DVDD:12391 0.0574016
rDVDD/2365 DVDD:12387 DVDD:12390 0.02916
rDVDD/2366 DVDD:12387 DVDD:12388 1.5
rDVDD/2367 DVDD:12385 DVDD:14493 0.0100984
rDVDD/2368 DVDD:12385 DVDD:12388 0.0574016
rDVDD/2369 DVDD:12384 DVDD:12387 0.02916
rDVDD/2370 DVDD:12384 DVDD:12385 1.5
rDVDD/2371 DVDD:12382 DVDD:14489 0.0186024
rDVDD/2372 DVDD:12382 DVDD:14493 0.0473032
rDVDD/2373 DVDD:12381 DVDD:12384 0.02916
rDVDD/2374 DVDD:12381 DVDD:12382 1.5
rDVDD/2375 DVDD:12379 DVDD:14485 0.0490748
rDVDD/2376 DVDD:12379 DVDD:14489 0.0387992
rDVDD/2377 DVDD:12378 DVDD:12381 0.02916
rDVDD/2378 DVDD:12378 DVDD:12379 1.5
rDVDD/2379 DVDD:12376 DVDD:14481 0.0575787
rDVDD/2380 DVDD:12376 DVDD:14485 0.00832677
rDVDD/2381 DVDD:12375 DVDD:12378 0.02916
rDVDD/2382 DVDD:12375 DVDD:12376 1.5
rDVDD/2383 DVDD:12368 DVDD:14474 0.00938976
rDVDD/2384 DVDD:12368 DVDD:14478 0.0565157
rDVDD/2385 DVDD:12367 DVDD:12368 2.25
rDVDD/2386 DVDD:12365 DVDD:14474 0.028878
rDVDD/2387 DVDD:12364 DVDD:12367 0.01944
rDVDD/2388 DVDD:12364 DVDD:12365 1.5
rDVDD/2389 DVDD:12362 DVDD:14469 0.00159449
rDVDD/2390 DVDD:12362 DVDD:12365 0.0574016
rDVDD/2391 DVDD:12361 DVDD:12364 0.02916
rDVDD/2392 DVDD:12361 DVDD:12362 1.5
rDVDD/2393 DVDD:12359 DVDD:14465 0.0497835
rDVDD/2394 DVDD:12359 DVDD:14469 0.0558071
rDVDD/2395 DVDD:12358 DVDD:12361 0.02916
rDVDD/2396 DVDD:12358 DVDD:12359 1.5
rDVDD/2397 DVDD:12356 DVDD:14465 0.00761811
rDVDD/2398 DVDD:12355 DVDD:12358 0.02916
rDVDD/2399 DVDD:12355 DVDD:12356 1.5
rDVDD/2400 DVDD:12353 DVDD:14460 0.0228543
rDVDD/2401 DVDD:12353 DVDD:12356 0.0574016
rDVDD/2402 DVDD:12352 DVDD:12355 0.02916
rDVDD/2403 DVDD:12352 DVDD:12353 1.5
rDVDD/2404 DVDD:12350 DVDD:14456 0.0313583
rDVDD/2405 DVDD:12350 DVDD:14460 0.0345472
rDVDD/2406 DVDD:12349 DVDD:12352 0.02916
rDVDD/2407 DVDD:12349 DVDD:12350 1.5
rDVDD/2408 DVDD:12347 DVDD:14456 0.0260433
rDVDD/2409 DVDD:12346 DVDD:12349 0.02916
rDVDD/2410 DVDD:12346 DVDD:12347 1.5
rDVDD/2411 DVDD:12344 DVDD:14451 0.00442913
rDVDD/2412 DVDD:12344 DVDD:12347 0.0574016
rDVDD/2413 DVDD:12343 DVDD:12346 0.02916
rDVDD/2414 DVDD:12343 DVDD:12344 1.5
rDVDD/2415 DVDD:12341 DVDD:14447 0.0129331
rDVDD/2416 DVDD:12341 DVDD:14451 0.0529724
rDVDD/2417 DVDD:12340 DVDD:12343 0.02916
rDVDD/2418 DVDD:12340 DVDD:12341 1.5
rDVDD/2419 DVDD:12328 DVDD:15007 0.0389764
rDVDD/2420 DVDD:12328 DVDD:12331 0.642857
rDVDD/2421 DVDD:12328 DVDD:15011 0.0885827
rDVDD/2422 DVDD:12327 DVDD:12328 0.5625
rDVDD/2423 DVDD:12315 DVDD:14722 0.0389764
rDVDD/2424 DVDD:12315 DVDD:12318 0.642857
rDVDD/2425 DVDD:12315 DVDD:14726 0.0666142
rDVDD/2426 DVDD:12314 DVDD:12315 0.5625
rDVDD/2427 DVDD:12301 DVDD:14437 0.0389764
rDVDD/2428 DVDD:12301 DVDD:12304 0.642857
rDVDD/2429 DVDD:12301 DVDD:14441 0.0666142
rDVDD/2430 DVDD:12300 DVDD:12301 0.5625
rDVDD/2431 DVDD:12288 DVDD:14158 0.0389764
rDVDD/2432 DVDD:12288 DVDD:12291 0.642857
rDVDD/2433 DVDD:12288 DVDD:14162 0.0885827
rDVDD/2434 DVDD:12287 DVDD:12288 0.5625
rDVDD/2435 DVDD:12275 DVDD:14968 0.051378
rDVDD/2436 DVDD:12275 DVDD:12278 0.642857
rDVDD/2437 DVDD:12275 DVDD:14972 0.0364961
rDVDD/2438 DVDD:12274 DVDD:12275 0.5625
rDVDD/2439 DVDD:12262 DVDD:14683 0.0733465
rDVDD/2440 DVDD:12262 DVDD:12265 0.642857
rDVDD/2441 DVDD:12262 DVDD:14687 0.0145276
rDVDD/2442 DVDD:12261 DVDD:12262 0.5625
rDVDD/2443 DVDD:12248 DVDD:14398 0.0733465
rDVDD/2444 DVDD:12248 DVDD:12251 0.642857
rDVDD/2445 DVDD:12248 DVDD:14402 0.0145276
rDVDD/2446 DVDD:12247 DVDD:12248 0.5625
rDVDD/2447 DVDD:12235 DVDD:14119 0.051378
rDVDD/2448 DVDD:12235 DVDD:12238 0.642857
rDVDD/2449 DVDD:12235 DVDD:14123 0.0364961
rDVDD/2450 DVDD:12234 DVDD:12235 0.5625
rDVDD/2451 DVDD:12224 DVDD:12226 2.28827
rDVDD/2452 DVDD:12223 DVDD:12226 0.01944
rDVDD/2453 DVDD:12223 DVDD:12224 1.5
rDVDD/2454 DVDD:12221 DVDD:12224 0.0574016
rDVDD/2455 DVDD:12220 DVDD:12223 0.02916
rDVDD/2456 DVDD:12220 DVDD:12221 1.5
rDVDD/2457 DVDD:12218 DVDD:14362 0.0210827
rDVDD/2458 DVDD:12218 DVDD:12221 0.0574016
rDVDD/2459 DVDD:12217 DVDD:12220 0.02916
rDVDD/2460 DVDD:12217 DVDD:12218 1.5
rDVDD/2461 DVDD:12215 DVDD:14358 0.0295866
rDVDD/2462 DVDD:12215 DVDD:14362 0.0363189
rDVDD/2463 DVDD:12214 DVDD:12217 0.02916
rDVDD/2464 DVDD:12214 DVDD:12215 1.5
rDVDD/2465 DVDD:12212 DVDD:14358 0.027815
rDVDD/2466 DVDD:12211 DVDD:12214 0.02916
rDVDD/2467 DVDD:12211 DVDD:12212 1.5
rDVDD/2468 DVDD:12209 DVDD:14353 0.00265748
rDVDD/2469 DVDD:12209 DVDD:12212 0.0574016
rDVDD/2470 DVDD:12208 DVDD:12211 0.02916
rDVDD/2471 DVDD:12208 DVDD:12209 1.5
rDVDD/2472 DVDD:12206 DVDD:14353 0.0547441
rDVDD/2473 DVDD:12205 DVDD:12208 0.02916
rDVDD/2474 DVDD:12205 DVDD:12206 1.5
rDVDD/2475 DVDD:12203 DVDD:12206 0.0574016
rDVDD/2476 DVDD:12202 DVDD:12205 0.02916
rDVDD/2477 DVDD:12202 DVDD:12203 1.5
rDVDD/2478 DVDD:12200 DVDD:12203 0.0574016
rDVDD/2479 DVDD:12199 DVDD:12202 0.02916
rDVDD/2480 DVDD:12199 DVDD:12200 1.5
rDVDD/2481 DVDD:12192 DVDD:12200 0.201969
rDVDD/2482 DVDD:12191 DVDD:12192 2.25
rDVDD/2483 DVDD:12189 DVDD:12192 0.0382677
rDVDD/2484 DVDD:12188 DVDD:12191 0.01944
rDVDD/2485 DVDD:12188 DVDD:12189 1.5
rDVDD/2486 DVDD:12186 DVDD:12189 0.0574016
rDVDD/2487 DVDD:12185 DVDD:12188 0.02916
rDVDD/2488 DVDD:12185 DVDD:12186 1.5
rDVDD/2489 DVDD:12183 DVDD:12186 0.0574016
rDVDD/2490 DVDD:12182 DVDD:12185 0.02916
rDVDD/2491 DVDD:12182 DVDD:12183 1.5
rDVDD/2492 DVDD:12180 DVDD:12183 0.0574016
rDVDD/2493 DVDD:12179 DVDD:12182 0.02916
rDVDD/2494 DVDD:12179 DVDD:12180 1.5
rDVDD/2495 DVDD:12177 DVDD:12180 0.0574016
rDVDD/2496 DVDD:12176 DVDD:12179 0.02916
rDVDD/2497 DVDD:12176 DVDD:12177 1.5
rDVDD/2498 DVDD:12174 DVDD:12177 0.0574016
rDVDD/2499 DVDD:12173 DVDD:12176 0.02916
rDVDD/2500 DVDD:12173 DVDD:12174 1.5
rDVDD/2501 DVDD:12171 DVDD:12174 0.0574016
rDVDD/2502 DVDD:12170 DVDD:12173 0.02916
rDVDD/2503 DVDD:12170 DVDD:12171 1.5
rDVDD/2504 DVDD:12168 DVDD:12171 0.0574016
rDVDD/2505 DVDD:12167 DVDD:12170 0.02916
rDVDD/2506 DVDD:12167 DVDD:12168 1.5
rDVDD/2507 DVDD:12165 DVDD:12168 0.0574016
rDVDD/2508 DVDD:12164 DVDD:12167 0.02916
rDVDD/2509 DVDD:12164 DVDD:12165 1.5
rDVDD/2510 DVDD:12157 DVDD:12165 0.201969
rDVDD/2511 DVDD:12156 DVDD:12157 2.25
rDVDD/2512 DVDD:12154 DVDD:12157 0.0382677
rDVDD/2513 DVDD:12153 DVDD:12156 0.01944
rDVDD/2514 DVDD:12153 DVDD:12154 1.5
rDVDD/2515 DVDD:12151 DVDD:12154 0.0574016
rDVDD/2516 DVDD:12150 DVDD:12153 0.02916
rDVDD/2517 DVDD:12150 DVDD:12151 1.5
rDVDD/2518 DVDD:12148 DVDD:14333 0.0395079
rDVDD/2519 DVDD:12148 DVDD:12151 0.0574016
rDVDD/2520 DVDD:12147 DVDD:12150 0.02916
rDVDD/2521 DVDD:12147 DVDD:12148 1.5
rDVDD/2522 DVDD:12145 DVDD:14329 0.0480118
rDVDD/2523 DVDD:12145 DVDD:14333 0.0178937
rDVDD/2524 DVDD:12144 DVDD:12147 0.02916
rDVDD/2525 DVDD:12144 DVDD:12145 1.5
rDVDD/2526 DVDD:12142 DVDD:14329 0.00938976
rDVDD/2527 DVDD:12141 DVDD:12144 0.02916
rDVDD/2528 DVDD:12141 DVDD:12142 1.5
rDVDD/2529 DVDD:12139 DVDD:14324 0.0210827
rDVDD/2530 DVDD:12139 DVDD:12142 0.0574016
rDVDD/2531 DVDD:12138 DVDD:12141 0.02916
rDVDD/2532 DVDD:12138 DVDD:12139 1.5
rDVDD/2533 DVDD:12136 DVDD:14324 0.0363189
rDVDD/2534 DVDD:12135 DVDD:12138 0.02916
rDVDD/2535 DVDD:12135 DVDD:12136 1.5
rDVDD/2536 DVDD:12133 DVDD:12136 0.0574016
rDVDD/2537 DVDD:12132 DVDD:12135 0.02916
rDVDD/2538 DVDD:12132 DVDD:12133 1.5
rDVDD/2539 DVDD:12130 DVDD:12133 0.0574016
rDVDD/2540 DVDD:12129 DVDD:12132 0.02916
rDVDD/2541 DVDD:12129 DVDD:12130 1.5
rDVDD/2542 DVDD:12122 DVDD:14317 0.016122
rDVDD/2543 DVDD:12122 DVDD:12130 0.201969
rDVDD/2544 DVDD:12121 DVDD:12122 2.25
rDVDD/2545 DVDD:12119 DVDD:14313 0.0437598
rDVDD/2546 DVDD:12119 DVDD:14317 0.0221457
rDVDD/2547 DVDD:12118 DVDD:12121 0.01944
rDVDD/2548 DVDD:12118 DVDD:12119 1.5
rDVDD/2549 DVDD:12116 DVDD:14313 0.0136417
rDVDD/2550 DVDD:12115 DVDD:12118 0.02916
rDVDD/2551 DVDD:12115 DVDD:12116 1.5
rDVDD/2552 DVDD:12113 DVDD:14308 0.0168307
rDVDD/2553 DVDD:12113 DVDD:12116 0.0574016
rDVDD/2554 DVDD:12112 DVDD:12115 0.02916
rDVDD/2555 DVDD:12112 DVDD:12113 1.5
rDVDD/2556 DVDD:12110 DVDD:14308 0.0405709
rDVDD/2557 DVDD:12109 DVDD:12112 0.02916
rDVDD/2558 DVDD:12109 DVDD:12110 1.5
rDVDD/2559 DVDD:12107 DVDD:14303 0.0317126
rDVDD/2560 DVDD:12107 DVDD:12110 0.0574016
rDVDD/2561 DVDD:12106 DVDD:12109 0.02916
rDVDD/2562 DVDD:12106 DVDD:12107 1.5
rDVDD/2563 DVDD:12104 DVDD:14303 0.025689
rDVDD/2564 DVDD:12103 DVDD:12106 0.02916
rDVDD/2565 DVDD:12103 DVDD:12104 1.5
rDVDD/2566 DVDD:12101 DVDD:14298 0.00478346
rDVDD/2567 DVDD:12101 DVDD:12104 0.0574016
rDVDD/2568 DVDD:12100 DVDD:12103 0.02916
rDVDD/2569 DVDD:12100 DVDD:12101 1.5
rDVDD/2570 DVDD:12098 DVDD:14294 0.0132874
rDVDD/2571 DVDD:12098 DVDD:14298 0.0526181
rDVDD/2572 DVDD:12097 DVDD:12100 0.02916
rDVDD/2573 DVDD:12097 DVDD:12098 1.5
rDVDD/2574 DVDD:12095 DVDD:14290 0.0855709
rDVDD/2575 DVDD:12095 DVDD:14294 0.0441142
rDVDD/2576 DVDD:12094 DVDD:12097 0.02916
rDVDD/2577 DVDD:12094 DVDD:12095 1.5
rDVDD/2578 DVDD:12087 DVDD:14284 0.00655512
rDVDD/2579 DVDD:12086 DVDD:12087 2.25
rDVDD/2580 DVDD:12084 DVDD:14279 0.0430512
rDVDD/2581 DVDD:12084 DVDD:12087 0.0382677
rDVDD/2582 DVDD:12083 DVDD:12086 0.01944
rDVDD/2583 DVDD:12083 DVDD:12084 1.5
rDVDD/2584 DVDD:12081 DVDD:14279 0.0143504
rDVDD/2585 DVDD:12080 DVDD:12083 0.02916
rDVDD/2586 DVDD:12080 DVDD:12081 1.5
rDVDD/2587 DVDD:12078 DVDD:12081 0.0574016
rDVDD/2588 DVDD:12077 DVDD:12080 0.02916
rDVDD/2589 DVDD:12077 DVDD:12078 1.5
rDVDD/2590 DVDD:12075 DVDD:12078 0.0574016
rDVDD/2591 DVDD:12074 DVDD:12077 0.02916
rDVDD/2592 DVDD:12074 DVDD:12075 1.5
rDVDD/2593 DVDD:12072 DVDD:12075 0.0574016
rDVDD/2594 DVDD:12071 DVDD:12074 0.02916
rDVDD/2595 DVDD:12071 DVDD:12072 1.5
rDVDD/2596 DVDD:12069 DVDD:12072 0.0574016
rDVDD/2597 DVDD:12068 DVDD:12071 0.02916
rDVDD/2598 DVDD:12068 DVDD:12069 1.5
rDVDD/2599 DVDD:12066 DVDD:12069 0.0574016
rDVDD/2600 DVDD:12065 DVDD:12068 0.02916
rDVDD/2601 DVDD:12065 DVDD:12066 1.5
rDVDD/2602 DVDD:12063 DVDD:12066 0.0574016
rDVDD/2603 DVDD:12062 DVDD:12065 0.02916
rDVDD/2604 DVDD:12062 DVDD:12063 1.5
rDVDD/2605 DVDD:12060 DVDD:12063 0.0574016
rDVDD/2606 DVDD:12059 DVDD:12062 0.02916
rDVDD/2607 DVDD:12059 DVDD:12060 1.5
rDVDD/2608 DVDD:12052 DVDD:12060 0.201969
rDVDD/2609 DVDD:12051 DVDD:12052 2.25
rDVDD/2610 DVDD:12049 DVDD:12052 0.0382677
rDVDD/2611 DVDD:12048 DVDD:12051 0.01944
rDVDD/2612 DVDD:12048 DVDD:12049 1.5
rDVDD/2613 DVDD:12046 DVDD:12049 0.0574016
rDVDD/2614 DVDD:12045 DVDD:12048 0.02916
rDVDD/2615 DVDD:12045 DVDD:12046 1.5
rDVDD/2616 DVDD:12043 DVDD:12046 0.0574016
rDVDD/2617 DVDD:12042 DVDD:12045 0.02916
rDVDD/2618 DVDD:12042 DVDD:12043 1.5
rDVDD/2619 DVDD:12040 DVDD:12043 0.0574016
rDVDD/2620 DVDD:12039 DVDD:12042 0.02916
rDVDD/2621 DVDD:12039 DVDD:12040 1.5
rDVDD/2622 DVDD:12037 DVDD:12040 0.0574016
rDVDD/2623 DVDD:12036 DVDD:12039 0.02916
rDVDD/2624 DVDD:12036 DVDD:12037 1.5
rDVDD/2625 DVDD:12034 DVDD:12037 0.0574016
rDVDD/2626 DVDD:12033 DVDD:12036 0.02916
rDVDD/2627 DVDD:12033 DVDD:12034 1.5
rDVDD/2628 DVDD:12031 DVDD:12034 0.0574016
rDVDD/2629 DVDD:12030 DVDD:12033 0.02916
rDVDD/2630 DVDD:12030 DVDD:12031 1.5
rDVDD/2631 DVDD:12028 DVDD:12031 0.0574016
rDVDD/2632 DVDD:12027 DVDD:12030 0.02916
rDVDD/2633 DVDD:12027 DVDD:12028 1.5
rDVDD/2634 DVDD:12025 DVDD:14258 0.14687
rDVDD/2635 DVDD:12025 DVDD:12028 0.0574016
rDVDD/2636 DVDD:12024 DVDD:12027 0.02916
rDVDD/2637 DVDD:12024 DVDD:12025 1.5
rDVDD/2638 DVDD:12017 DVDD:14254 0.0108071
rDVDD/2639 DVDD:12017 DVDD:14258 0.0550984
rDVDD/2640 DVDD:12016 DVDD:12017 2.25
rDVDD/2641 DVDD:12014 DVDD:14254 0.0274606
rDVDD/2642 DVDD:12013 DVDD:12016 0.01944
rDVDD/2643 DVDD:12013 DVDD:12014 1.5
rDVDD/2644 DVDD:12011 DVDD:14249 0.00301181
rDVDD/2645 DVDD:12011 DVDD:12014 0.0574016
rDVDD/2646 DVDD:12010 DVDD:12013 0.02916
rDVDD/2647 DVDD:12010 DVDD:12011 1.5
rDVDD/2648 DVDD:12008 DVDD:14245 0.0115157
rDVDD/2649 DVDD:12008 DVDD:14249 0.0543898
rDVDD/2650 DVDD:12007 DVDD:12010 0.02916
rDVDD/2651 DVDD:12007 DVDD:12008 1.5
rDVDD/2652 DVDD:12005 DVDD:14241 0.0419882
rDVDD/2653 DVDD:12005 DVDD:14245 0.0458858
rDVDD/2654 DVDD:12004 DVDD:12007 0.02916
rDVDD/2655 DVDD:12004 DVDD:12005 1.5
rDVDD/2656 DVDD:12002 DVDD:14241 0.0154134
rDVDD/2657 DVDD:12001 DVDD:12004 0.02916
rDVDD/2658 DVDD:12001 DVDD:12002 1.5
rDVDD/2659 DVDD:11999 DVDD:14236 0.0150591
rDVDD/2660 DVDD:11999 DVDD:12002 0.0574016
rDVDD/2661 DVDD:11998 DVDD:12001 0.02916
rDVDD/2662 DVDD:11998 DVDD:11999 1.5
rDVDD/2663 DVDD:11996 DVDD:14236 0.0423425
rDVDD/2664 DVDD:11995 DVDD:11998 0.02916
rDVDD/2665 DVDD:11995 DVDD:11996 1.5
rDVDD/2666 DVDD:11993 DVDD:14231 0.028878
rDVDD/2667 DVDD:11993 DVDD:11996 0.0574016
rDVDD/2668 DVDD:11992 DVDD:11995 0.02916
rDVDD/2669 DVDD:11992 DVDD:11993 1.5
rDVDD/2670 DVDD:11990 DVDD:14227 0.0154134
rDVDD/2671 DVDD:11990 DVDD:14231 0.0285236
rDVDD/2672 DVDD:11989 DVDD:11992 0.02916
rDVDD/2673 DVDD:11989 DVDD:11990 1.5
rDVDD/2674 DVDD:11982 DVDD:14221 0.0327756
rDVDD/2675 DVDD:11981 DVDD:11982 2.25
rDVDD/2676 DVDD:11979 DVDD:11982 0.0382677
rDVDD/2677 DVDD:11978 DVDD:11981 0.01944
rDVDD/2678 DVDD:11978 DVDD:11979 1.5
rDVDD/2679 DVDD:11976 DVDD:11979 0.0574016
rDVDD/2680 DVDD:11975 DVDD:11978 0.02916
rDVDD/2681 DVDD:11975 DVDD:11976 1.5
rDVDD/2682 DVDD:11973 DVDD:11976 0.0574016
rDVDD/2683 DVDD:11972 DVDD:11975 0.02916
rDVDD/2684 DVDD:11972 DVDD:11973 1.5
rDVDD/2685 DVDD:11970 DVDD:11973 0.0574016
rDVDD/2686 DVDD:11969 DVDD:11972 0.02916
rDVDD/2687 DVDD:11969 DVDD:11970 1.5
rDVDD/2688 DVDD:11967 DVDD:11970 0.0574016
rDVDD/2689 DVDD:11966 DVDD:11969 0.02916
rDVDD/2690 DVDD:11966 DVDD:11967 1.5
rDVDD/2691 DVDD:11964 DVDD:14211 0.0540354
rDVDD/2692 DVDD:11964 DVDD:11967 0.0574016
rDVDD/2693 DVDD:11963 DVDD:11966 0.02916
rDVDD/2694 DVDD:11963 DVDD:11964 1.5
rDVDD/2695 DVDD:11961 DVDD:14211 0.00336614
rDVDD/2696 DVDD:11960 DVDD:11963 0.02916
rDVDD/2697 DVDD:11960 DVDD:11961 1.5
rDVDD/2698 DVDD:11958 DVDD:14206 0.0051378
rDVDD/2699 DVDD:11958 DVDD:11961 0.0574016
rDVDD/2700 DVDD:11957 DVDD:11960 0.02916
rDVDD/2701 DVDD:11957 DVDD:11958 1.5
rDVDD/2702 DVDD:11955 DVDD:14202 0.0356102
rDVDD/2703 DVDD:11955 DVDD:14206 0.0522638
rDVDD/2704 DVDD:11954 DVDD:11957 0.02916
rDVDD/2705 DVDD:11954 DVDD:11955 1.5
rDVDD/2706 DVDD:11947 DVDD:14196 0.0125787
rDVDD/2707 DVDD:11946 DVDD:11947 2.25
rDVDD/2708 DVDD:11944 DVDD:14191 0.0370276
rDVDD/2709 DVDD:11944 DVDD:11947 0.0382677
rDVDD/2710 DVDD:11943 DVDD:11946 0.01944
rDVDD/2711 DVDD:11943 DVDD:11944 1.5
rDVDD/2712 DVDD:11941 DVDD:14191 0.020374
rDVDD/2713 DVDD:11940 DVDD:11943 0.02916
rDVDD/2714 DVDD:11940 DVDD:11941 1.5
rDVDD/2715 DVDD:11938 DVDD:14186 0.0497835
rDVDD/2716 DVDD:11938 DVDD:11941 0.0574016
rDVDD/2717 DVDD:11937 DVDD:11940 0.02916
rDVDD/2718 DVDD:11937 DVDD:11938 1.5
rDVDD/2719 DVDD:11935 DVDD:14182 0.0363189
rDVDD/2720 DVDD:11935 DVDD:14186 0.00761811
rDVDD/2721 DVDD:11934 DVDD:11937 0.02916
rDVDD/2722 DVDD:11934 DVDD:11935 1.5
rDVDD/2723 DVDD:11932 DVDD:14178 0.0448228
rDVDD/2724 DVDD:11932 DVDD:14182 0.0210827
rDVDD/2725 DVDD:11931 DVDD:11934 0.02916
rDVDD/2726 DVDD:11931 DVDD:11932 1.5
rDVDD/2727 DVDD:11929 DVDD:14178 0.0125787
rDVDD/2728 DVDD:11928 DVDD:11931 0.02916
rDVDD/2729 DVDD:11928 DVDD:11929 1.5
rDVDD/2730 DVDD:11926 DVDD:14173 0.0178937
rDVDD/2731 DVDD:11926 DVDD:11929 0.0574016
rDVDD/2732 DVDD:11925 DVDD:11928 0.02916
rDVDD/2733 DVDD:11925 DVDD:11926 1.5
rDVDD/2734 DVDD:11923 DVDD:14169 0.0263976
rDVDD/2735 DVDD:11923 DVDD:14173 0.0395079
rDVDD/2736 DVDD:11922 DVDD:11925 0.02916
rDVDD/2737 DVDD:11922 DVDD:11923 1.5
rDVDD/2738 DVDD:11920 DVDD:14165 0.0568701
rDVDD/2739 DVDD:11920 DVDD:14169 0.0310039
rDVDD/2740 DVDD:11919 DVDD:11922 0.02916
rDVDD/2741 DVDD:11919 DVDD:11920 1.5
rDVDD/2742 DVDD:11907 DVDD:11910 0.0486
rDVDD/2743 DVDD:11903 DVDD:11910 4.5
rDVDD/2744 DVDD:11903 DVDD:15001 0.00797244
rDVDD/2745 DVDD:11902 DVDD:11903 1.5
rDVDD/2746 DVDD:11900 DVDD:14996 0.0607677
rDVDD/2747 DVDD:11900 DVDD:11907 1.5
rDVDD/2748 DVDD:11900 DVDD:11903 0.0191339
rDVDD/2749 DVDD:11899 DVDD:11902 0.0486
rDVDD/2750 DVDD:11899 DVDD:11900 1.5
rDVDD/2751 DVDD:11881 DVDD:11884 0.0486
rDVDD/2752 DVDD:11879 DVDD:11884 4.5
rDVDD/2753 DVDD:11879 DVDD:14719 0.0299409
rDVDD/2754 DVDD:11878 DVDD:11881 0.0972
rDVDD/2755 DVDD:11878 DVDD:11879 1.5
rDVDD/2756 DVDD:11876 DVDD:14714 0.0387992
rDVDD/2757 DVDD:11876 DVDD:11881 1.5
rDVDD/2758 DVDD:11876 DVDD:11879 0.0191339
rDVDD/2759 DVDD:11875 DVDD:11878 0.0486
rDVDD/2760 DVDD:11875 DVDD:11876 1.5
rDVDD/2761 DVDD:11853 DVDD:14434 0.0299409
rDVDD/2762 DVDD:11852 DVDD:11853 1.5
rDVDD/2763 DVDD:11850 DVDD:14429 0.0387992
rDVDD/2764 DVDD:11850 DVDD:11853 0.0191339
rDVDD/2765 DVDD:11849 DVDD:11852 0.0486
rDVDD/2766 DVDD:11849 DVDD:11850 1.5
rDVDD/2767 DVDD:11831 DVDD:11834 0.0486
rDVDD/2768 DVDD:11827 DVDD:11834 4.5
rDVDD/2769 DVDD:11827 DVDD:14152 0.00797244
rDVDD/2770 DVDD:11826 DVDD:11827 1.5
rDVDD/2771 DVDD:11824 DVDD:14147 0.0607677
rDVDD/2772 DVDD:11824 DVDD:11831 1.5
rDVDD/2773 DVDD:11824 DVDD:11827 0.0191339
rDVDD/2774 DVDD:11823 DVDD:11826 0.0486
rDVDD/2775 DVDD:11823 DVDD:11824 1.5
rDVDD/2776 DVDD:11811 DVDD:11814 0.0486
rDVDD/2777 DVDD:11807 DVDD:11814 4.5
rDVDD/2778 DVDD:11807 DVDD:14993 0.0086811
rDVDD/2779 DVDD:11806 DVDD:11807 1.5
rDVDD/2780 DVDD:11804 DVDD:14988 0.0600591
rDVDD/2781 DVDD:11804 DVDD:11811 1.5
rDVDD/2782 DVDD:11804 DVDD:11807 0.0191339
rDVDD/2783 DVDD:11803 DVDD:11806 0.0486
rDVDD/2784 DVDD:11803 DVDD:11804 1.5
rDVDD/2785 DVDD:11785 DVDD:11788 0.0486
rDVDD/2786 DVDD:11783 DVDD:11788 4.5
rDVDD/2787 DVDD:11783 DVDD:14711 0.0306496
rDVDD/2788 DVDD:11782 DVDD:11785 0.0972
rDVDD/2789 DVDD:11782 DVDD:11783 1.5
rDVDD/2790 DVDD:11780 DVDD:14706 0.0380905
rDVDD/2791 DVDD:11780 DVDD:11785 1.5
rDVDD/2792 DVDD:11780 DVDD:11783 0.0191339
rDVDD/2793 DVDD:11779 DVDD:11782 0.0486
rDVDD/2794 DVDD:11779 DVDD:11780 1.5
rDVDD/2795 DVDD:11757 DVDD:14426 0.0306496
rDVDD/2796 DVDD:11756 DVDD:11757 1.5
rDVDD/2797 DVDD:11754 DVDD:14421 0.0380905
rDVDD/2798 DVDD:11754 DVDD:11757 0.0191339
rDVDD/2799 DVDD:11753 DVDD:11756 0.0486
rDVDD/2800 DVDD:11753 DVDD:11754 1.5
rDVDD/2801 DVDD:11735 DVDD:11738 0.0486
rDVDD/2802 DVDD:11731 DVDD:11738 4.5
rDVDD/2803 DVDD:11731 DVDD:14144 0.0086811
rDVDD/2804 DVDD:11730 DVDD:11731 1.5
rDVDD/2805 DVDD:11728 DVDD:14139 0.0600591
rDVDD/2806 DVDD:11728 DVDD:11735 1.5
rDVDD/2807 DVDD:11728 DVDD:11731 0.0191339
rDVDD/2808 DVDD:11727 DVDD:11730 0.0486
rDVDD/2809 DVDD:11727 DVDD:11728 1.5
rDVDD/2810 DVDD:11715 DVDD:11718 0.0486
rDVDD/2811 DVDD:11711 DVDD:14984 0.0125787
rDVDD/2812 DVDD:11711 DVDD:11718 4.5
rDVDD/2813 DVDD:11711 DVDD:14988 0.0752953
rDVDD/2814 DVDD:11710 DVDD:11711 1.5
rDVDD/2815 DVDD:11708 DVDD:14980 0.121004
rDVDD/2816 DVDD:11708 DVDD:11715 1.5
rDVDD/2817 DVDD:11708 DVDD:14984 0.00655512
rDVDD/2818 DVDD:11707 DVDD:11710 0.0486
rDVDD/2819 DVDD:11707 DVDD:11708 1.5
rDVDD/2820 DVDD:11689 DVDD:11692 0.0486
rDVDD/2821 DVDD:11687 DVDD:11692 4.5
rDVDD/2822 DVDD:11687 DVDD:14703 0.0313583
rDVDD/2823 DVDD:11686 DVDD:11689 0.0972
rDVDD/2824 DVDD:11686 DVDD:11687 1.5
rDVDD/2825 DVDD:11684 DVDD:14698 0.0373819
rDVDD/2826 DVDD:11684 DVDD:11689 1.5
rDVDD/2827 DVDD:11684 DVDD:11687 0.0191339
rDVDD/2828 DVDD:11683 DVDD:11686 0.0486
rDVDD/2829 DVDD:11683 DVDD:11684 1.5
rDVDD/2830 DVDD:11661 DVDD:14418 0.0313583
rDVDD/2831 DVDD:11660 DVDD:11661 1.5
rDVDD/2832 DVDD:11658 DVDD:14413 0.0373819
rDVDD/2833 DVDD:11658 DVDD:11661 0.0191339
rDVDD/2834 DVDD:11657 DVDD:11660 0.0486
rDVDD/2835 DVDD:11657 DVDD:11658 1.5
rDVDD/2836 DVDD:11639 DVDD:11642 0.0486
rDVDD/2837 DVDD:11635 DVDD:14135 0.0125787
rDVDD/2838 DVDD:11635 DVDD:11642 4.5
rDVDD/2839 DVDD:11635 DVDD:14139 0.0752953
rDVDD/2840 DVDD:11634 DVDD:11635 1.5
rDVDD/2841 DVDD:11632 DVDD:14131 0.121004
rDVDD/2842 DVDD:11632 DVDD:11639 1.5
rDVDD/2843 DVDD:11632 DVDD:14135 0.00655512
rDVDD/2844 DVDD:11631 DVDD:11634 0.0486
rDVDD/2845 DVDD:11631 DVDD:11632 1.5
rDVDD/2846 DVDD:11619 DVDD:11622 0.0486
rDVDD/2847 DVDD:11615 DVDD:11622 4.5
rDVDD/2848 DVDD:11615 DVDD:14980 0.0143504
rDVDD/2849 DVDD:11614 DVDD:11615 1.5
rDVDD/2850 DVDD:11612 DVDD:14975 0.0543898
rDVDD/2851 DVDD:11612 DVDD:11619 1.5
rDVDD/2852 DVDD:11612 DVDD:11615 0.0191339
rDVDD/2853 DVDD:11611 DVDD:11614 0.0486
rDVDD/2854 DVDD:11611 DVDD:11612 1.5
rDVDD/2855 DVDD:11593 DVDD:11596 0.0486
rDVDD/2856 DVDD:11591 DVDD:11596 4.5
rDVDD/2857 DVDD:11591 DVDD:14695 0.0143504
rDVDD/2858 DVDD:11590 DVDD:11593 0.0972
rDVDD/2859 DVDD:11590 DVDD:11591 1.5
rDVDD/2860 DVDD:11588 DVDD:14690 0.0763583
rDVDD/2861 DVDD:11588 DVDD:11593 1.5
rDVDD/2862 DVDD:11588 DVDD:11591 0.0191339
rDVDD/2863 DVDD:11587 DVDD:11590 0.0486
rDVDD/2864 DVDD:11587 DVDD:11588 1.5
rDVDD/2865 DVDD:11565 DVDD:14410 0.0143504
rDVDD/2866 DVDD:11564 DVDD:11565 1.5
rDVDD/2867 DVDD:11562 DVDD:14405 0.0763583
rDVDD/2868 DVDD:11562 DVDD:11565 0.0191339
rDVDD/2869 DVDD:11561 DVDD:11564 0.0486
rDVDD/2870 DVDD:11561 DVDD:11562 1.5
rDVDD/2871 DVDD:11543 DVDD:11546 0.0486
rDVDD/2872 DVDD:11539 DVDD:11546 4.5
rDVDD/2873 DVDD:11539 DVDD:14131 0.0143504
rDVDD/2874 DVDD:11538 DVDD:11539 1.5
rDVDD/2875 DVDD:11536 DVDD:14126 0.0543898
rDVDD/2876 DVDD:11536 DVDD:11543 1.5
rDVDD/2877 DVDD:11536 DVDD:11539 0.0191339
rDVDD/2878 DVDD:11535 DVDD:11538 0.0486
rDVDD/2879 DVDD:11535 DVDD:11536 1.5
rDVDD/2880 DVDD:11527 DVDD:11528 4.5
rDVDD/2881 DVDD:11525 DVDD:11528 0.0558
rDVDD/2882 DVDD:11524 DVDD:11527 0.01116
rDVDD/2883 DVDD:11524 DVDD:11525 1.5
rDVDD/2884 DVDD:11522 DVDD:11525 0.0558
rDVDD/2885 DVDD:11521 DVDD:11524 0.01116
rDVDD/2886 DVDD:11521 DVDD:11522 1.5
rDVDD/2887 DVDD:11519 DVDD:11522 0.1116
rDVDD/2888 DVDD:11518 DVDD:11521 0.02232
rDVDD/2889 DVDD:11518 DVDD:11519 1.5
rDVDD/2890 DVDD:11516 DVDD:11519 0.0558
rDVDD/2891 DVDD:11515 DVDD:11518 0.01116
rDVDD/2892 DVDD:11515 DVDD:11516 1.5
rDVDD/2893 DVDD:11513 DVDD:11516 0.1116
rDVDD/2894 DVDD:11512 DVDD:11515 0.02232
rDVDD/2895 DVDD:11512 DVDD:11513 1.5
rDVDD/2896 DVDD:11510 DVDD:11513 0.0558
rDVDD/2897 DVDD:11509 DVDD:11512 0.01116
rDVDD/2898 DVDD:11509 DVDD:11510 1.5
rDVDD/2899 DVDD:11507 DVDD:11510 0.1116
rDVDD/2900 DVDD:11506 DVDD:11509 0.02232
rDVDD/2901 DVDD:11506 DVDD:11507 1.5
rDVDD/2902 DVDD:11504 DVDD:11507 0.0558
rDVDD/2903 DVDD:11503 DVDD:11506 0.01116
rDVDD/2904 DVDD:11503 DVDD:11504 1.5
rDVDD/2905 DVDD:11501 DVDD:11504 0.1116
rDVDD/2906 DVDD:11500 DVDD:11503 0.02232
rDVDD/2907 DVDD:11500 DVDD:11501 1.5
rDVDD/2908 DVDD:11498 DVDD:11501 0.0558
rDVDD/2909 DVDD:11497 DVDD:11500 0.01116
rDVDD/2910 DVDD:11497 DVDD:11498 1.5
rDVDD/2911 DVDD:11495 DVDD:11498 0.1116
rDVDD/2912 DVDD:11494 DVDD:11497 0.02232
rDVDD/2913 DVDD:11494 DVDD:11495 1.5
rDVDD/2914 DVDD:11492 DVDD:11495 0.0558
rDVDD/2915 DVDD:11491 DVDD:11494 0.01116
rDVDD/2916 DVDD:11491 DVDD:11492 1.5
rDVDD/2917 DVDD:11489 DVDD:11492 0.1116
rDVDD/2918 DVDD:11488 DVDD:11491 0.02232
rDVDD/2919 DVDD:11488 DVDD:11489 1.5
rDVDD/2920 DVDD:11486 DVDD:11489 0.0558
rDVDD/2921 DVDD:11485 DVDD:11488 0.01116
rDVDD/2922 DVDD:11485 DVDD:11486 1.5
rDVDD/2923 DVDD:11483 DVDD:11486 0.1116
rDVDD/2924 DVDD:11482 DVDD:11485 0.02232
rDVDD/2925 DVDD:11482 DVDD:11483 1.5
rDVDD/2926 DVDD:11480 DVDD:11483 0.0558
rDVDD/2927 DVDD:11479 DVDD:11482 0.01116
rDVDD/2928 DVDD:11479 DVDD:11480 1.5
rDVDD/2929 DVDD:11477 DVDD:11480 0.1116
rDVDD/2930 DVDD:11476 DVDD:11479 0.02232
rDVDD/2931 DVDD:11476 DVDD:11477 1.5
rDVDD/2932 DVDD:11469 DVDD:11477 0.3816
rDVDD/2933 DVDD:11468 DVDD:11469 4.5
rDVDD/2934 DVDD:11466 DVDD:11469 0.0558
rDVDD/2935 DVDD:11465 DVDD:11468 0.01116
rDVDD/2936 DVDD:11465 DVDD:11466 1.5
rDVDD/2937 DVDD:11463 DVDD:11466 0.0558
rDVDD/2938 DVDD:11462 DVDD:11465 0.01116
rDVDD/2939 DVDD:11462 DVDD:11463 1.5
rDVDD/2940 DVDD:11460 DVDD:11463 0.1116
rDVDD/2941 DVDD:11459 DVDD:11462 0.02232
rDVDD/2942 DVDD:11459 DVDD:11460 1.5
rDVDD/2943 DVDD:11457 DVDD:11460 0.0558
rDVDD/2944 DVDD:11456 DVDD:11459 0.01116
rDVDD/2945 DVDD:11456 DVDD:11457 1.5
rDVDD/2946 DVDD:11454 DVDD:13858 0.05265
rDVDD/2947 DVDD:11454 DVDD:11457 0.1116
rDVDD/2948 DVDD:11453 DVDD:11456 0.02232
rDVDD/2949 DVDD:11453 DVDD:11454 1.5
rDVDD/2950 DVDD:11451 DVDD:13854 0.05265
rDVDD/2951 DVDD:11451 DVDD:13858 0.00315
rDVDD/2952 DVDD:11450 DVDD:11453 0.01116
rDVDD/2953 DVDD:11450 DVDD:11451 1.5
rDVDD/2954 DVDD:11448 DVDD:13854 0.05895
rDVDD/2955 DVDD:11448 DVDD:13834 1.5
rDVDD/2956 DVDD:11447 DVDD:11450 0.02232
rDVDD/2957 DVDD:11447 DVDD:11448 1.5
rDVDD/2958 DVDD:11445 DVDD:13847 0.05265
rDVDD/2959 DVDD:11445 DVDD:11448 0.0558
rDVDD/2960 DVDD:11444 DVDD:11447 0.01116
rDVDD/2961 DVDD:11444 DVDD:11445 1.5
rDVDD/2962 DVDD:11442 DVDD:13847 0.05895
rDVDD/2963 DVDD:11442 DVDD:13834 1.5
rDVDD/2964 DVDD:11441 DVDD:11444 0.02232
rDVDD/2965 DVDD:11441 DVDD:11442 1.5
rDVDD/2966 DVDD:11439 DVDD:13840 0.05265
rDVDD/2967 DVDD:11439 DVDD:11442 0.0558
rDVDD/2968 DVDD:11438 DVDD:11441 0.01116
rDVDD/2969 DVDD:11438 DVDD:11439 1.5
rDVDD/2970 DVDD:11436 DVDD:13840 0.05895
rDVDD/2971 DVDD:11436 DVDD:13834 1.5
rDVDD/2972 DVDD:11435 DVDD:11438 0.02232
rDVDD/2973 DVDD:11435 DVDD:11436 1.5
rDVDD/2974 DVDD:11433 DVDD:13833 0.05265
rDVDD/2975 DVDD:11433 DVDD:11436 0.0558
rDVDD/2976 DVDD:11432 DVDD:11435 0.01116
rDVDD/2977 DVDD:11432 DVDD:11433 1.5
rDVDD/2978 DVDD:11430 DVDD:13833 0.05895
rDVDD/2979 DVDD:11429 DVDD:11432 0.02232
rDVDD/2980 DVDD:11429 DVDD:11430 1.5
rDVDD/2981 DVDD:11427 DVDD:11430 0.0558
rDVDD/2982 DVDD:11426 DVDD:11429 0.01116
rDVDD/2983 DVDD:11426 DVDD:11427 1.5
rDVDD/2984 DVDD:11424 DVDD:11427 0.1116
rDVDD/2985 DVDD:11423 DVDD:11426 0.02232
rDVDD/2986 DVDD:11423 DVDD:11424 1.5
rDVDD/2987 DVDD:11421 DVDD:11424 0.0558
rDVDD/2988 DVDD:11420 DVDD:11423 0.01116
rDVDD/2989 DVDD:11420 DVDD:11421 1.5
rDVDD/2990 DVDD:11418 DVDD:11421 0.1116
rDVDD/2991 DVDD:11417 DVDD:11420 0.02232
rDVDD/2992 DVDD:11417 DVDD:11418 1.5
rDVDD/2993 DVDD:11410 DVDD:11418 0.3816
rDVDD/2994 DVDD:11409 DVDD:11410 4.5
rDVDD/2995 DVDD:11407 DVDD:11410 0.0558
rDVDD/2996 DVDD:11406 DVDD:11409 0.01116
rDVDD/2997 DVDD:11406 DVDD:11407 1.5
rDVDD/2998 DVDD:11404 DVDD:11407 0.0558
rDVDD/2999 DVDD:11404 DVDD:13753 1.5
rDVDD/3000 DVDD:11403 DVDD:11406 0.01116
rDVDD/3001 DVDD:11403 DVDD:11404 1.5
rDVDD/3002 DVDD:11401 DVDD:11404 0.1116
rDVDD/3003 DVDD:11401 DVDD:13753 1.5
rDVDD/3004 DVDD:11400 DVDD:11403 0.02232
rDVDD/3005 DVDD:11400 DVDD:11401 1.5
rDVDD/3006 DVDD:11398 DVDD:11401 0.0558
rDVDD/3007 DVDD:11398 DVDD:13753 1.5
rDVDD/3008 DVDD:11397 DVDD:11400 0.01116
rDVDD/3009 DVDD:11397 DVDD:11398 1.5
rDVDD/3010 DVDD:11395 DVDD:11398 0.1116
rDVDD/3011 DVDD:11395 DVDD:13753 1.5
rDVDD/3012 DVDD:11394 DVDD:11397 0.02232
rDVDD/3013 DVDD:11394 DVDD:11395 1.5
rDVDD/3014 DVDD:11392 DVDD:11395 0.0558
rDVDD/3015 DVDD:11392 DVDD:13753 1.5
rDVDD/3016 DVDD:11391 DVDD:11394 0.01116
rDVDD/3017 DVDD:11391 DVDD:11392 1.5
rDVDD/3018 DVDD:11389 DVDD:11392 0.1116
rDVDD/3019 DVDD:11389 DVDD:13753 1.5
rDVDD/3020 DVDD:11388 DVDD:11391 0.02232
rDVDD/3021 DVDD:11388 DVDD:11389 1.5
rDVDD/3022 DVDD:11386 DVDD:11389 0.0558
rDVDD/3023 DVDD:11386 DVDD:13753 1.5
rDVDD/3024 DVDD:11385 DVDD:11388 0.01116
rDVDD/3025 DVDD:11385 DVDD:11386 1.5
rDVDD/3026 DVDD:11383 DVDD:11386 0.1116
rDVDD/3027 DVDD:11382 DVDD:11385 0.02232
rDVDD/3028 DVDD:11382 DVDD:11383 1.5
rDVDD/3029 DVDD:11380 DVDD:13800 0.04545
rDVDD/3030 DVDD:11380 DVDD:11383 0.0558
rDVDD/3031 DVDD:11379 DVDD:11382 0.01116
rDVDD/3032 DVDD:11379 DVDD:11380 1.5
rDVDD/3033 DVDD:11377 DVDD:13800 0.06615
rDVDD/3034 DVDD:11377 DVDD:13753 1.5
rDVDD/3035 DVDD:11376 DVDD:11379 0.02232
rDVDD/3036 DVDD:11376 DVDD:11377 1.5
rDVDD/3037 DVDD:11374 DVDD:13793 0.04545
rDVDD/3038 DVDD:11374 DVDD:11377 0.0558
rDVDD/3039 DVDD:11373 DVDD:11376 0.01116
rDVDD/3040 DVDD:11373 DVDD:11374 1.5
rDVDD/3041 DVDD:11371 DVDD:13793 0.06615
rDVDD/3042 DVDD:11371 DVDD:13753 1.5
rDVDD/3043 DVDD:11370 DVDD:11373 0.02232
rDVDD/3044 DVDD:11370 DVDD:11371 1.5
rDVDD/3045 DVDD:11368 DVDD:13786 0.04545
rDVDD/3046 DVDD:11368 DVDD:11371 0.0558
rDVDD/3047 DVDD:11367 DVDD:11370 0.01116
rDVDD/3048 DVDD:11367 DVDD:11368 1.5
rDVDD/3049 DVDD:11365 DVDD:13786 0.06615
rDVDD/3050 DVDD:11365 DVDD:13753 1.5
rDVDD/3051 DVDD:11364 DVDD:11367 0.02232
rDVDD/3052 DVDD:11364 DVDD:11365 1.5
rDVDD/3053 DVDD:11362 DVDD:13779 0.04545
rDVDD/3054 DVDD:11362 DVDD:11365 0.0558
rDVDD/3055 DVDD:11361 DVDD:11364 0.01116
rDVDD/3056 DVDD:11361 DVDD:11362 1.5
rDVDD/3057 DVDD:11359 DVDD:13773 0.20745
rDVDD/3058 DVDD:11359 DVDD:13779 0.06615
rDVDD/3059 DVDD:11359 DVDD:13753 1.5
rDVDD/3060 DVDD:11358 DVDD:11361 0.02232
rDVDD/3061 DVDD:11358 DVDD:11359 1.5
rDVDD/3062 DVDD:11351 DVDD:13767 0.00675
rDVDD/3063 DVDD:11350 DVDD:11351 4.5
rDVDD/3064 DVDD:11348 DVDD:11351 0.0558
rDVDD/3065 DVDD:11348 DVDD:13753 1.5
rDVDD/3066 DVDD:11347 DVDD:11350 0.01116
rDVDD/3067 DVDD:11347 DVDD:11348 1.5
rDVDD/3068 DVDD:11345 DVDD:13759 0.04905
rDVDD/3069 DVDD:11345 DVDD:11348 0.0558
rDVDD/3070 DVDD:11344 DVDD:11347 0.01116
rDVDD/3071 DVDD:11344 DVDD:11345 1.5
rDVDD/3072 DVDD:11342 DVDD:13759 0.06255
rDVDD/3073 DVDD:11342 DVDD:13753 1.5
rDVDD/3074 DVDD:11341 DVDD:11344 0.02232
rDVDD/3075 DVDD:11341 DVDD:11342 1.5
rDVDD/3076 DVDD:11339 DVDD:13752 0.04905
rDVDD/3077 DVDD:11339 DVDD:11342 0.0558
rDVDD/3078 DVDD:11338 DVDD:11341 0.01116
rDVDD/3079 DVDD:11338 DVDD:11339 1.5
rDVDD/3080 DVDD:11336 DVDD:13752 0.06255
rDVDD/3081 DVDD:11335 DVDD:11338 0.02232
rDVDD/3082 DVDD:11335 DVDD:11336 1.5
rDVDD/3083 DVDD:11333 DVDD:11336 0.0558
rDVDD/3084 DVDD:11332 DVDD:11335 0.01116
rDVDD/3085 DVDD:11332 DVDD:11333 1.5
rDVDD/3086 DVDD:11330 DVDD:11333 0.1116
rDVDD/3087 DVDD:11329 DVDD:11332 0.02232
rDVDD/3088 DVDD:11329 DVDD:11330 1.5
rDVDD/3089 DVDD:11327 DVDD:11330 0.0558
rDVDD/3090 DVDD:11326 DVDD:11329 0.01116
rDVDD/3091 DVDD:11326 DVDD:11327 1.5
rDVDD/3092 DVDD:11324 DVDD:11327 0.1116
rDVDD/3093 DVDD:11323 DVDD:11326 0.02232
rDVDD/3094 DVDD:11323 DVDD:11324 1.5
rDVDD/3095 DVDD:11321 DVDD:11324 0.0558
rDVDD/3096 DVDD:11320 DVDD:11323 0.01116
rDVDD/3097 DVDD:11320 DVDD:11321 1.5
rDVDD/3098 DVDD:11318 DVDD:11321 0.1116
rDVDD/3099 DVDD:11317 DVDD:11320 0.02232
rDVDD/3100 DVDD:11317 DVDD:11318 1.5
rDVDD/3101 DVDD:11315 DVDD:11318 0.0558
rDVDD/3102 DVDD:11314 DVDD:11317 0.01116
rDVDD/3103 DVDD:11314 DVDD:11315 1.5
rDVDD/3104 DVDD:11312 DVDD:11315 0.1116
rDVDD/3105 DVDD:11311 DVDD:11314 0.02232
rDVDD/3106 DVDD:11311 DVDD:11312 1.5
rDVDD/3107 DVDD:11309 DVDD:11312 0.0558
rDVDD/3108 DVDD:11308 DVDD:11311 0.01116
rDVDD/3109 DVDD:11308 DVDD:11309 1.5
rDVDD/3110 DVDD:11306 DVDD:11309 0.1116
rDVDD/3111 DVDD:11305 DVDD:11308 0.02232
rDVDD/3112 DVDD:11305 DVDD:11306 1.5
rDVDD/3113 DVDD:11303 DVDD:11306 0.0558
rDVDD/3114 DVDD:11302 DVDD:11305 0.01116
rDVDD/3115 DVDD:11302 DVDD:11303 1.5
rDVDD/3116 DVDD:11300 DVDD:11303 0.1116
rDVDD/3117 DVDD:11299 DVDD:11302 0.02232
rDVDD/3118 DVDD:11299 DVDD:11300 1.5
rDVDD/3119 DVDD:11289 DVDD:15743 0.00261161
rDVDD/3120 DVDD:11289 DVDD:15749 0.0222991
rDVDD/3121 DVDD:11288 DVDD:11289 1.5
rDVDD/3122 DVDD:11286 DVDD:13735 0.0275223
rDVDD/3123 DVDD:11286 DVDD:15743 0.0472098
rDVDD/3124 DVDD:11285 DVDD:11288 0.02232
rDVDD/3125 DVDD:11285 DVDD:11286 0.5625
rDVDD/3126 DVDD:11283 DVDD:13731 0.0275223
rDVDD/3127 DVDD:11283 DVDD:13735 0.0472098
rDVDD/3128 DVDD:11282 DVDD:11285 0.03348
rDVDD/3129 DVDD:11282 DVDD:11283 0.5625
rDVDD/3130 DVDD:11280 DVDD:15740 0.0275223
rDVDD/3131 DVDD:11280 DVDD:13731 0.0222991
rDVDD/3132 DVDD:11279 DVDD:11282 0.02232
rDVDD/3133 DVDD:11279 DVDD:11280 0.5625
rDVDD/3134 DVDD:11277 DVDD:15733 0.00261161
rDVDD/3135 DVDD:11277 DVDD:15740 0.0222991
rDVDD/3136 DVDD:11276 DVDD:11279 0.02232
rDVDD/3137 DVDD:11276 DVDD:11277 1.5
rDVDD/3138 DVDD:11249 DVDD:13725 0.0310669
rDVDD/3139 DVDD:11248 DVDD:11249 4.5
rDVDD/3140 DVDD:11246 DVDD:13720 0.0156276
rDVDD/3141 DVDD:11246 DVDD:11249 0.0233473
rDVDD/3142 DVDD:11245 DVDD:11248 0.01116
rDVDD/3143 DVDD:11245 DVDD:11246 0.5625
rDVDD/3144 DVDD:11243 DVDD:13716 0.0389749
rDVDD/3145 DVDD:11243 DVDD:13720 0.0544142
rDVDD/3146 DVDD:11242 DVDD:11245 0.03348
rDVDD/3147 DVDD:11242 DVDD:11243 0.5625
rDVDD/3148 DVDD:11240 DVDD:13712 0.0389749
rDVDD/3149 DVDD:11240 DVDD:13716 0.0310669
rDVDD/3150 DVDD:11239 DVDD:11242 0.03348
rDVDD/3151 DVDD:11239 DVDD:11240 0.5625
rDVDD/3152 DVDD:11237 DVDD:13712 0.00771967
rDVDD/3153 DVDD:11236 DVDD:11239 0.02232
rDVDD/3154 DVDD:11236 DVDD:11237 0.5625
rDVDD/3155 DVDD:11234 DVDD:13707 0.0156276
rDVDD/3156 DVDD:11234 DVDD:11237 0.0700418
rDVDD/3157 DVDD:11233 DVDD:11236 0.03348
rDVDD/3158 DVDD:11233 DVDD:11234 0.5625
rDVDD/3159 DVDD:11231 DVDD:13703 0.0389749
rDVDD/3160 DVDD:11231 DVDD:13707 0.0544142
rDVDD/3161 DVDD:11230 DVDD:11233 0.03348
rDVDD/3162 DVDD:11230 DVDD:11231 0.5625
rDVDD/3163 DVDD:11228 DVDD:13703 0.00771967
rDVDD/3164 DVDD:11227 DVDD:11230 0.02232
rDVDD/3165 DVDD:11227 DVDD:11228 0.5625
rDVDD/3166 DVDD:11223 DVDD:13698 0.0589331
rDVDD/3167 DVDD:11223 DVDD:15768 0.0344561
rDVDD/3168 DVDD:11222 DVDD:11223 0.5
rDVDD/3169 DVDD:11215 DVDD:15714 0.0160042
rDVDD/3170 DVDD:11215 DVDD:15721 0.0073431
rDVDD/3171 DVDD:11214 DVDD:11215 1.5
rDVDD/3172 DVDD:11206 DVDD:15704 0.0103556
rDVDD/3173 DVDD:11206 DVDD:15710 0.0129916
rDVDD/3174 DVDD:11205 DVDD:11206 1.5
rDVDD/3175 DVDD:11203 DVDD:13686 0.0570502
rDVDD/3176 DVDD:11203 DVDD:13690 0.0129916
rDVDD/3177 DVDD:11202 DVDD:11205 0.02232
rDVDD/3178 DVDD:11202 DVDD:11203 0.5625
rDVDD/3179 DVDD:11200 DVDD:13686 0.0129916
rDVDD/3180 DVDD:11199 DVDD:11202 0.03348
rDVDD/3181 DVDD:11199 DVDD:11200 0.5625
rDVDD/3182 DVDD:11197 DVDD:13681 0.0337029
rDVDD/3183 DVDD:11197 DVDD:11200 0.0466946
rDVDD/3184 DVDD:11196 DVDD:11199 0.02232
rDVDD/3185 DVDD:11196 DVDD:11197 0.5625
rDVDD/3186 DVDD:11189 DVDD:13675 0.00922594
rDVDD/3187 DVDD:11188 DVDD:11189 0.9
rDVDD/3188 DVDD:11186 DVDD:13670 0.0374686
rDVDD/3189 DVDD:11186 DVDD:11189 0.0466946
rDVDD/3190 DVDD:11185 DVDD:11188 0.02232
rDVDD/3191 DVDD:11185 DVDD:11186 0.5625
rDVDD/3192 DVDD:11183 DVDD:13670 0.00922594
rDVDD/3193 DVDD:11182 DVDD:11185 0.02232
rDVDD/3194 DVDD:11182 DVDD:11183 0.5625
rDVDD/3195 DVDD:11178 DVDD:15763 0.0137448
rDVDD/3196 DVDD:11177 DVDD:11178 1.5
rDVDD/3197 DVDD:11175 DVDD:13665 0.00960251
rDVDD/3198 DVDD:11175 DVDD:11178 0.0233473
rDVDD/3199 DVDD:11174 DVDD:11177 0.01116
rDVDD/3200 DVDD:11174 DVDD:11175 2.25
rDVDD/3201 DVDD:11172 DVDD:13661 0.0329498
rDVDD/3202 DVDD:11172 DVDD:13665 0.037092
rDVDD/3203 DVDD:11171 DVDD:11174 0.02232
rDVDD/3204 DVDD:11171 DVDD:11172 0.5625
rDVDD/3205 DVDD:11169 DVDD:13661 0.0137448
rDVDD/3206 DVDD:11168 DVDD:11171 0.02232
rDVDD/3207 DVDD:11168 DVDD:11169 0.5625
rDVDD/3208 DVDD:11166 DVDD:13656 0.00960251
rDVDD/3209 DVDD:11166 DVDD:11169 0.0700418
rDVDD/3210 DVDD:11165 DVDD:11168 0.03348
rDVDD/3211 DVDD:11165 DVDD:11166 0.5625
rDVDD/3212 DVDD:11163 DVDD:13652 0.00960251
rDVDD/3213 DVDD:11163 DVDD:13656 0.0604393
rDVDD/3214 DVDD:11162 DVDD:11165 0.03348
rDVDD/3215 DVDD:11162 DVDD:11163 0.5625
rDVDD/3216 DVDD:11160 DVDD:13648 0.0562971
rDVDD/3217 DVDD:11160 DVDD:13652 0.037092
rDVDD/3218 DVDD:11159 DVDD:11162 0.02232
rDVDD/3219 DVDD:11159 DVDD:11160 0.5625
rDVDD/3220 DVDD:11149 DVDD:16209 0.0627189
rDVDD/3221 DVDD:11149 DVDD:16206 0.0576923
rDVDD/3222 DVDD:11144 DVDD:11149 0.00376991
rDVDD/3223 DVDD:11144 DVDD:16200 0.0112876
rDVDD/3224 DVDD:11141 DVDD:11144 0.0201062
rDVDD/3225 DVDD:11141 DVDD:16195 0.0140333
rDVDD/3226 DVDD:11137 DVDD:16188 0.00701663
rDVDD/3227 DVDD:11137 DVDD:16195 0.0452389
rDVDD/3228 DVDD:11136 DVDD:11141 0.0201062
rDVDD/3229 DVDD:11136 DVDD:11137 0.00701663
rDVDD/3230 DVDD:11134 DVDD:16183 0.0140333
rDVDD/3231 DVDD:11134 DVDD:16177 0.0452389
rDVDD/3232 DVDD:11134 DVDD:11137 0.0452389
rDVDD/3233 DVDD:11133 DVDD:11136 0.0201062
rDVDD/3234 DVDD:11133 DVDD:11134 0.0140333
rDVDD/3235 DVDD:11128 DVDD:11133 0.0201062
rDVDD/3236 DVDD:11128 DVDD:16177 0.00701663
rDVDD/3237 DVDD:11126 DVDD 0.0333717
rDVDD/3238 DVDD:11126 DVDD:16172 0.0140333
rDVDD/3239 DVDD:11126 DVDD:16177 0.0452389
rDVDD/3240 DVDD:11125 DVDD:11128 0.0201062
rDVDD/3241 DVDD:11125 DVDD:11126 0.0140333
rDVDD/3242 DVDD DVDD:11125 0.0148319
rDVDD/3243 DVDD DVDD:16163 0.0193076
rDVDD/3244 DVDD:11112 DVDD:16160 0.0581321
rDVDD/3245 DVDD:11112 DVDD:16157 0.0531496
rDVDD/3246 DVDD:11107 DVDD:11112 0.00498246
rDVDD/3247 DVDD:11107 DVDD:16151 0.0108521
rDVDD/3248 DVDD:11104 DVDD:11107 0.0199298
rDVDD/3249 DVDD:11104 DVDD:16147 0.0136364
rDVDD/3250 DVDD:11100 DVDD:16140 0.00681818
rDVDD/3251 DVDD:11100 DVDD:16147 0.0448421
rDVDD/3252 DVDD:11099 DVDD:11104 0.0199298
rDVDD/3253 DVDD:11099 DVDD:11100 0.00681818
rDVDD/3254 DVDD:11097 DVDD:16136 0.0136364
rDVDD/3255 DVDD:11097 DVDD:16131 0.0448421
rDVDD/3256 DVDD:11097 DVDD:11100 0.0448421
rDVDD/3257 DVDD:11096 DVDD:11099 0.0199298
rDVDD/3258 DVDD:11096 DVDD:11097 0.0136364
rDVDD/3259 DVDD:11091 DVDD:11096 0.0199298
rDVDD/3260 DVDD:11091 DVDD:16131 0.00681818
rDVDD/3261 DVDD:11089 DVDD 0.0302763
rDVDD/3262 DVDD:11089 DVDD:16126 0.0136364
rDVDD/3263 DVDD:11089 DVDD:16131 0.0448421
rDVDD/3264 DVDD:11088 DVDD:11091 0.0199298
rDVDD/3265 DVDD:11088 DVDD:11089 0.0136364
rDVDD/3266 DVDD DVDD:11088 0.0134561
rDVDD/3267 DVDD DVDD:16117 0.0188644
rDVDD/3268 DVDD:11080 DVDD 0.00874739
rDVDD/3269 DVDD:11080 DVDD:15436 0.00823043
rDVDD/3270 DVDD DVDD:11080 0.00543306
rDVDD/3272 DVDD:11073 DVDD 0.00843845
rDVDD/3273 DVDD:11073 DVDD:16106 0.00154533
rDVDD/3274 DVDD:11073 DVDD 0.0104254
rDVDD/3275 DVDD:11072 DVDD 0.00463351
rDVDD/3276 DVDD:11072 DVDD:11073 0.00154533
rDVDD/3277 DVDD DVDD:11072 0.00375042
rDVDD/3279 DVDD:11066 DVDD 0.00584341
rDVDD/3280 DVDD:11066 DVDD 0.0086747
rDVDD/3281 DVDD:11066 DVDD 0.00540075
rDVDD/3282 DVDD:11060 DVDD:16083 0.166179
rDVDD/3283 DVDD:11060 DVDD:16084 0.0456429
rDVDD/3284 DVDD:11056 DVDD:11060 0.140821
rDVDD/3285 DVDD:11056 DVDD:16084 0.143617
rDVDD/3286 DVDD:11053 DVDD:11056 0.0162286
rDVDD/3287 DVDD:11053 DVDD:16080 0.143617
rDVDD/3288 DVDD:11050 DVDD:11053 0.00405714
rDVDD/3289 DVDD:11050 DVDD:16077 0.143617
rDVDD/3290 DVDD:11047 DVDD:11050 0.0202857
rDVDD/3291 DVDD:11047 DVDD:16073 0.143617
rDVDD/3292 DVDD:11042 DVDD:11047 0.0162286
rDVDD/3293 DVDD:11042 DVDD:16068 0.0718085
rDVDD/3294 DVDD:11039 DVDD:11042 0.0202857
rDVDD/3295 DVDD:11039 DVDD:16065 0.143617
rDVDD/3296 DVDD:11035 DVDD:16058 0.0718085
rDVDD/3297 DVDD:11035 DVDD:16065 0.0365143
rDVDD/3298 DVDD:11034 DVDD:11039 0.0162286
rDVDD/3299 DVDD:11034 DVDD:11035 0.0718085
rDVDD/3300 DVDD:11032 DVDD:16055 0.143617
rDVDD/3301 DVDD:11032 DVDD:11035 0.0456429
rDVDD/3302 DVDD:11031 DVDD:11034 0.0202857
rDVDD/3303 DVDD:11031 DVDD:11032 0.143617
rDVDD/3304 DVDD:11027 DVDD:16050 0.0718085
rDVDD/3305 DVDD:11027 DVDD:11032 0.0456429
rDVDD/3306 DVDD:11026 DVDD:11031 0.0202857
rDVDD/3307 DVDD:11026 DVDD:11027 0.0718085
rDVDD/3308 DVDD:11024 DVDD:16046 0.143617
rDVDD/3309 DVDD:11024 DVDD:11027 0.0456429
rDVDD/3310 DVDD:11023 DVDD:11026 0.0202857
rDVDD/3311 DVDD:11023 DVDD:11024 0.143617
rDVDD/3312 DVDD:11019 DVDD:16041 0.0718085
rDVDD/3313 DVDD:11019 DVDD:11024 0.0365143
rDVDD/3314 DVDD:11018 DVDD:11023 0.0162286
rDVDD/3315 DVDD:11018 DVDD:11019 0.0718085
rDVDD/3316 DVDD:11016 DVDD:16038 0.143617
rDVDD/3317 DVDD:11016 DVDD:11019 0.0456429
rDVDD/3318 DVDD:11015 DVDD:11018 0.0202857
rDVDD/3319 DVDD:11015 DVDD:11016 0.143617
rDVDD/3320 DVDD:11013 DVDD:16035 0.143617
rDVDD/3321 DVDD:11013 DVDD:11016 0.0365143
rDVDD/3322 DVDD:11012 DVDD:11015 0.0162286
rDVDD/3323 DVDD:11012 DVDD:11013 0.143617
rDVDD/3324 DVDD:11010 DVDD:16032 0.143617
rDVDD/3325 DVDD:11010 DVDD:11013 0.00912857
rDVDD/3326 DVDD:11009 DVDD:11012 0.00405714
rDVDD/3327 DVDD:11009 DVDD:11010 0.143617
rDVDD/3328 DVDD:11007 DVDD:16028 0.143617
rDVDD/3329 DVDD:11007 DVDD:16024 0.0365143
rDVDD/3330 DVDD:11007 DVDD:11010 0.0456429
rDVDD/3331 DVDD:11006 DVDD:11009 0.0202857
rDVDD/3332 DVDD:11006 DVDD:11007 0.143617
rDVDD/3333 DVDD:11001 DVDD:11006 0.0162286
rDVDD/3334 DVDD:11001 DVDD:16024 0.0718085
rDVDD/3335 DVDD:10998 DVDD:11001 0.0202857
rDVDD/3336 DVDD:10998 DVDD:16021 0.143617
rDVDD/3337 DVDD:10994 DVDD:16015 0.0718085
rDVDD/3338 DVDD:10994 DVDD:16021 0.0365143
rDVDD/3339 DVDD:10993 DVDD:10998 0.0162286
rDVDD/3340 DVDD:10993 DVDD:10994 0.0718085
rDVDD/3341 DVDD:10991 DVDD:16011 0.143617
rDVDD/3342 DVDD:10991 DVDD:10994 0.0456429
rDVDD/3343 DVDD:10990 DVDD:10993 0.0202857
rDVDD/3344 DVDD:10990 DVDD:10991 0.143617
rDVDD/3345 DVDD:10986 DVDD:16006 0.0718085
rDVDD/3346 DVDD:10986 DVDD:16003 0.0456429
rDVDD/3347 DVDD:10986 DVDD:10991 0.0456429
rDVDD/3348 DVDD:10985 DVDD:10990 0.0202857
rDVDD/3349 DVDD:10985 DVDD:10986 0.0718085
rDVDD/3350 DVDD:10982 DVDD:10985 0.0202857
rDVDD/3351 DVDD:10982 DVDD:16003 0.143617
rDVDD/3352 DVDD:10977 DVDD:10982 0.0162286
rDVDD/3353 DVDD:10977 DVDD:15998 0.0718085
rDVDD/3354 DVDD DVDD:10977 0.0194857
rDVDD/3355 DVDD:10972 DVDD 0.0008
rDVDD/3356 DVDD:10972 DVDD:15990 0.143617
rDVDD/3357 DVDD:10972 DVDD:15986 0.159846
rDVDD/3358 DVDD:10963 DVDD:15976 0.166179
rDVDD/3359 DVDD:10963 DVDD:15977 0.0456429
rDVDD/3360 DVDD:10959 DVDD:10963 0.140821
rDVDD/3361 DVDD:10959 DVDD:15977 0.143617
rDVDD/3362 DVDD:10956 DVDD:10959 0.0162286
rDVDD/3363 DVDD:10956 DVDD:15973 0.143617
rDVDD/3364 DVDD:10953 DVDD:10956 0.00405714
rDVDD/3365 DVDD:10953 DVDD:15970 0.143617
rDVDD/3366 DVDD:10950 DVDD:10953 0.0202857
rDVDD/3367 DVDD:10950 DVDD:15966 0.143617
rDVDD/3368 DVDD:10945 DVDD:10950 0.0162286
rDVDD/3369 DVDD:10945 DVDD:15961 0.0718085
rDVDD/3370 DVDD:10942 DVDD:10945 0.0202857
rDVDD/3371 DVDD:10942 DVDD:15958 0.143617
rDVDD/3372 DVDD:10938 DVDD:15951 0.0718085
rDVDD/3373 DVDD:10938 DVDD:15958 0.0365143
rDVDD/3374 DVDD:10937 DVDD:10942 0.0162286
rDVDD/3375 DVDD:10937 DVDD:10938 0.0718085
rDVDD/3376 DVDD:10935 DVDD:15948 0.143617
rDVDD/3377 DVDD:10935 DVDD:10938 0.0456429
rDVDD/3378 DVDD:10934 DVDD:10937 0.0202857
rDVDD/3379 DVDD:10934 DVDD:10935 0.143617
rDVDD/3380 DVDD:10930 DVDD:15943 0.0718085
rDVDD/3381 DVDD:10930 DVDD:10935 0.0456429
rDVDD/3382 DVDD:10929 DVDD:10934 0.0202857
rDVDD/3383 DVDD:10929 DVDD:10930 0.0718085
rDVDD/3384 DVDD:10927 DVDD:15939 0.143617
rDVDD/3385 DVDD:10927 DVDD:10930 0.0456429
rDVDD/3386 DVDD:10926 DVDD:10929 0.0202857
rDVDD/3387 DVDD:10926 DVDD:10927 0.143617
rDVDD/3388 DVDD:10922 DVDD:15934 0.0718085
rDVDD/3389 DVDD:10922 DVDD:10927 0.0365143
rDVDD/3390 DVDD:10921 DVDD:10926 0.0162286
rDVDD/3391 DVDD:10921 DVDD:10922 0.0718085
rDVDD/3392 DVDD:10919 DVDD:15931 0.143617
rDVDD/3393 DVDD:10919 DVDD:10922 0.0456429
rDVDD/3394 DVDD:10918 DVDD:10921 0.0202857
rDVDD/3395 DVDD:10918 DVDD:10919 0.143617
rDVDD/3396 DVDD:10916 DVDD:15928 0.143617
rDVDD/3397 DVDD:10916 DVDD:10919 0.0365143
rDVDD/3398 DVDD:10915 DVDD:10918 0.0162286
rDVDD/3399 DVDD:10915 DVDD:10916 0.143617
rDVDD/3400 DVDD:10913 DVDD:15925 0.143617
rDVDD/3401 DVDD:10913 DVDD:10916 0.00912857
rDVDD/3402 DVDD:10912 DVDD:10915 0.00405714
rDVDD/3403 DVDD:10912 DVDD:10913 0.143617
rDVDD/3404 DVDD:10910 DVDD:15921 0.143617
rDVDD/3405 DVDD:10910 DVDD:15917 0.0365143
rDVDD/3406 DVDD:10910 DVDD:10913 0.0456429
rDVDD/3407 DVDD:10909 DVDD:10912 0.0202857
rDVDD/3408 DVDD:10909 DVDD:10910 0.143617
rDVDD/3409 DVDD:10904 DVDD:10909 0.0162286
rDVDD/3410 DVDD:10904 DVDD:15917 0.0718085
rDVDD/3411 DVDD:10901 DVDD:10904 0.0202857
rDVDD/3412 DVDD:10901 DVDD:15914 0.143617
rDVDD/3413 DVDD:10897 DVDD:15908 0.0718085
rDVDD/3414 DVDD:10897 DVDD:15914 0.0365143
rDVDD/3415 DVDD:10896 DVDD:10901 0.0162286
rDVDD/3416 DVDD:10896 DVDD:10897 0.0718085
rDVDD/3417 DVDD:10894 DVDD:15904 0.143617
rDVDD/3418 DVDD:10894 DVDD:10897 0.0456429
rDVDD/3419 DVDD:10893 DVDD:10896 0.0202857
rDVDD/3420 DVDD:10893 DVDD:10894 0.143617
rDVDD/3421 DVDD:10889 DVDD:15899 0.0718085
rDVDD/3422 DVDD:10889 DVDD:15896 0.0456429
rDVDD/3423 DVDD:10889 DVDD:10894 0.0456429
rDVDD/3424 DVDD:10888 DVDD:10893 0.0202857
rDVDD/3425 DVDD:10888 DVDD:10889 0.0718085
rDVDD/3426 DVDD:10885 DVDD:10888 0.0202857
rDVDD/3427 DVDD:10885 DVDD:15896 0.143617
rDVDD/3428 DVDD:10880 DVDD:10885 0.0162286
rDVDD/3429 DVDD:10880 DVDD:15891 0.0718085
rDVDD/3430 DVDD DVDD:10880 0.0194857
rDVDD/3431 DVDD:10875 DVDD 0.0008
rDVDD/3432 DVDD:10875 DVDD:15884 0.143617
rDVDD/3433 DVDD:10875 DVDD:15880 0.159846
rDVDD/3434 DVDD:10866 DVDD:15870 0.166179
rDVDD/3435 DVDD:10866 DVDD:15871 0.0456429
rDVDD/3436 DVDD:10862 DVDD:10866 0.140821
rDVDD/3437 DVDD:10862 DVDD:15871 0.143617
rDVDD/3438 DVDD:10859 DVDD:10862 0.0162286
rDVDD/3439 DVDD:10859 DVDD:15867 0.143617
rDVDD/3440 DVDD:10856 DVDD:10859 0.00405714
rDVDD/3441 DVDD:10856 DVDD:15864 0.143617
rDVDD/3442 DVDD:10853 DVDD:10856 0.0202857
rDVDD/3443 DVDD:10853 DVDD:15860 0.143617
rDVDD/3444 DVDD:10848 DVDD:10853 0.0162286
rDVDD/3445 DVDD:10848 DVDD:15855 0.0718085
rDVDD/3446 DVDD:10845 DVDD:10848 0.0202857
rDVDD/3447 DVDD:10845 DVDD:15852 0.143617
rDVDD/3448 DVDD:10841 DVDD:15845 0.0718085
rDVDD/3449 DVDD:10841 DVDD:15852 0.0365143
rDVDD/3450 DVDD:10840 DVDD:10845 0.0162286
rDVDD/3451 DVDD:10840 DVDD:10841 0.0718085
rDVDD/3452 DVDD:10838 DVDD:15842 0.143617
rDVDD/3453 DVDD:10838 DVDD:10841 0.0456429
rDVDD/3454 DVDD:10837 DVDD:10840 0.0202857
rDVDD/3455 DVDD:10837 DVDD:10838 0.143617
rDVDD/3456 DVDD:10833 DVDD:15837 0.0718085
rDVDD/3457 DVDD:10833 DVDD:10838 0.0456429
rDVDD/3458 DVDD:10832 DVDD:10837 0.0202857
rDVDD/3459 DVDD:10832 DVDD:10833 0.0718085
rDVDD/3460 DVDD:10830 DVDD:15833 0.143617
rDVDD/3461 DVDD:10830 DVDD:10833 0.0456429
rDVDD/3462 DVDD:10829 DVDD:10832 0.0202857
rDVDD/3463 DVDD:10829 DVDD:10830 0.143617
rDVDD/3464 DVDD:10825 DVDD:15828 0.0718085
rDVDD/3465 DVDD:10825 DVDD:10830 0.0365143
rDVDD/3466 DVDD:10824 DVDD:10829 0.0162286
rDVDD/3467 DVDD:10824 DVDD:10825 0.0718085
rDVDD/3468 DVDD:10822 DVDD:15825 0.143617
rDVDD/3469 DVDD:10822 DVDD:10825 0.0456429
rDVDD/3470 DVDD:10821 DVDD:10824 0.0202857
rDVDD/3471 DVDD:10821 DVDD:10822 0.143617
rDVDD/3472 DVDD:10819 DVDD:15822 0.143617
rDVDD/3473 DVDD:10819 DVDD:10822 0.0365143
rDVDD/3474 DVDD:10818 DVDD:10821 0.0162286
rDVDD/3475 DVDD:10818 DVDD:10819 0.143617
rDVDD/3476 DVDD:10816 DVDD:15819 0.143617
rDVDD/3477 DVDD:10816 DVDD:10819 0.00912857
rDVDD/3478 DVDD:10815 DVDD:10818 0.00405714
rDVDD/3479 DVDD:10815 DVDD:10816 0.143617
rDVDD/3480 DVDD:10813 DVDD:15815 0.143617
rDVDD/3481 DVDD:10813 DVDD:15811 0.0365143
rDVDD/3482 DVDD:10813 DVDD:10816 0.0456429
rDVDD/3483 DVDD:10812 DVDD:10815 0.0202857
rDVDD/3484 DVDD:10812 DVDD:10813 0.143617
rDVDD/3485 DVDD:10807 DVDD:10812 0.0162286
rDVDD/3486 DVDD:10807 DVDD:15811 0.0718085
rDVDD/3487 DVDD:10804 DVDD:10807 0.0202857
rDVDD/3488 DVDD:10804 DVDD:15808 0.143617
rDVDD/3489 DVDD:10800 DVDD:15802 0.0718085
rDVDD/3490 DVDD:10800 DVDD:15808 0.0365143
rDVDD/3491 DVDD:10799 DVDD:10804 0.0162286
rDVDD/3492 DVDD:10799 DVDD:10800 0.0718085
rDVDD/3493 DVDD:10797 DVDD:15798 0.143617
rDVDD/3494 DVDD:10797 DVDD:10800 0.0456429
rDVDD/3495 DVDD:10796 DVDD:10799 0.0202857
rDVDD/3496 DVDD:10796 DVDD:10797 0.143617
rDVDD/3497 DVDD:10792 DVDD:15793 0.0718085
rDVDD/3498 DVDD:10792 DVDD:15790 0.0456429
rDVDD/3499 DVDD:10792 DVDD:10797 0.0456429
rDVDD/3500 DVDD:10791 DVDD:10796 0.0202857
rDVDD/3501 DVDD:10791 DVDD:10792 0.0718085
rDVDD/3502 DVDD:10788 DVDD:10791 0.0202857
rDVDD/3503 DVDD:10788 DVDD:15790 0.143617
rDVDD/3504 DVDD:10783 DVDD:10788 0.0162286
rDVDD/3505 DVDD:10783 DVDD:15785 0.0718085
rDVDD/3506 DVDD DVDD:10783 0.0194857
rDVDD/3507 DVDD:10778 DVDD 0.0008
rDVDD/3508 DVDD:10778 DVDD:15777 0.143617
rDVDD/3509 DVDD:10778 DVDD:15773 0.159846
rDVDD/3510 DVDD:10771 DVDD:10772 1.5
rDVDD/3511 DVDD:10771 DVDD:11528 0.371457
rDVDD/3512 DVDD:10766 DVDD:11300 0.392617
rDVDD/3513 DVDD:10766 DVDD:10767 1.5
rDVDD/3514 DVDD:10761 DVDD:15729 0.228015
rDVDD/3515 DVDD:10761 DVDD:10762 1.5
rDVDD/3516 DVDD:10758 DVDD:11227 0.02232
rDVDD/3517 DVDD:10757 DVDD:11228 0.0466946
rDVDD/3518 DVDD:10757 DVDD:10758 1.5
rDVDD/3519 DVDD:10753 DVDD:11182 0.02232
rDVDD/3520 DVDD:10752 DVDD:11183 0.0466946
rDVDD/3521 DVDD:10752 DVDD:10753 1.5
rDVDD/3522 DVDD:10731 DVDD:10734 0.03348
rDVDD/3523 DVDD:10730 DVDD:10734 0.665833
rDVDD/3524 DVDD:10730 DVDD:10731 0.5625
rDVDD/3525 DVDD:10728 DVDD:11288 0.02232
rDVDD/3526 DVDD:10728 DVDD:10731 0.02232
rDVDD/3527 DVDD:10727 DVDD:15749 0.0421811
rDVDD/3528 DVDD:10727 DVDD:10730 0.0688889
rDVDD/3529 DVDD:10727 DVDD:10728 0.5625
rDVDD/3530 DVDD:10724 DVDD:11276 0.02232
rDVDD/3531 DVDD:10723 DVDD:15733 0.0694033
rDVDD/3532 DVDD:10723 DVDD:10724 0.9
rDVDD/3533 DVDD:10721 DVDD:10724 0.02232
rDVDD/3534 DVDD:10720 DVDD:10723 0.0688889
rDVDD/3535 DVDD:10720 DVDD:10721 0.5625
rDVDD/3536 DVDD:10718 DVDD:10772 0.02232
rDVDD/3537 DVDD:10718 DVDD:10721 0.02232
rDVDD/3538 DVDD:10717 DVDD:10720 0.0688889
rDVDD/3539 DVDD:10717 DVDD:10718 0.5625
rDVDD/3540 DVDD:10717 DVDD:10771 0.0710706
rDVDD/3541 DVDD:10713 DVDD:10767 0.02232
rDVDD/3542 DVDD:10712 DVDD:10766 0.0603243
rDVDD/3543 DVDD:10712 DVDD:10713 0.5625
rDVDD/3544 DVDD:10710 DVDD:10713 0.03348
rDVDD/3545 DVDD:10709 DVDD:10712 0.0904865
rDVDD/3546 DVDD:10709 DVDD:10710 0.5625
rDVDD/3547 DVDD:10707 DVDD:10710 0.02232
rDVDD/3548 DVDD:10706 DVDD:10709 0.0603243
rDVDD/3549 DVDD:10706 DVDD:10707 0.5625
rDVDD/3550 DVDD:10704 DVDD:10707 0.03348
rDVDD/3551 DVDD:10703 DVDD:10706 0.0904865
rDVDD/3552 DVDD:10703 DVDD:10704 0.5625
rDVDD/3553 DVDD:10701 DVDD:10704 0.03348
rDVDD/3554 DVDD:10700 DVDD:10703 0.0904865
rDVDD/3555 DVDD:10700 DVDD:10701 0.5625
rDVDD/3556 DVDD:10698 DVDD:10701 0.02232
rDVDD/3557 DVDD:10697 DVDD:10700 0.0603243
rDVDD/3558 DVDD:10697 DVDD:10698 0.5625
rDVDD/3559 DVDD:10695 DVDD:10698 0.03348
rDVDD/3560 DVDD:10694 DVDD:10697 0.0904865
rDVDD/3561 DVDD:10694 DVDD:10695 0.5625
rDVDD/3562 DVDD:10692 DVDD:10695 0.03348
rDVDD/3563 DVDD:10691 DVDD:10694 0.0904865
rDVDD/3564 DVDD:10691 DVDD:10692 0.5625
rDVDD/3565 DVDD:10689 DVDD:10762 0.02232
rDVDD/3566 DVDD:10689 DVDD:10692 0.02232
rDVDD/3567 DVDD:10688 DVDD:10761 0.0603243
rDVDD/3568 DVDD:10688 DVDD:10691 0.0603243
rDVDD/3569 DVDD:10688 DVDD:10689 0.5625
rDVDD/3570 DVDD:10684 DVDD:11222 0.03348
rDVDD/3571 DVDD:10684 DVDD:10758 0.02232
rDVDD/3572 DVDD:10683 DVDD:15768 0.048715
rDVDD/3573 DVDD:10683 DVDD:10757 0.0585047
rDVDD/3574 DVDD:10683 DVDD:10684 0.5
rDVDD/3575 DVDD:10679 DVDD:11214 0.02232
rDVDD/3576 DVDD:10678 DVDD:15714 0.0423906
rDVDD/3577 DVDD:10678 DVDD:10679 0.5625
rDVDD/3578 DVDD:10676 DVDD:10679 0.03348
rDVDD/3579 DVDD:10675 DVDD:10678 0.0904865
rDVDD/3580 DVDD:10675 DVDD:10676 0.5625
rDVDD/3581 DVDD:10673 DVDD:10676 0.02232
rDVDD/3582 DVDD:10672 DVDD:10675 0.0603243
rDVDD/3583 DVDD:10672 DVDD:10673 0.5625
rDVDD/3584 DVDD:10670 DVDD:10673 0.03348
rDVDD/3585 DVDD:10669 DVDD:10672 0.0904865
rDVDD/3586 DVDD:10669 DVDD:10670 0.5625
rDVDD/3587 DVDD:10667 DVDD:10670 0.03348
rDVDD/3588 DVDD:10666 DVDD:10669 0.0904865
rDVDD/3589 DVDD:10666 DVDD:10667 0.5625
rDVDD/3590 DVDD:10664 DVDD:11205 0.02232
rDVDD/3591 DVDD:10664 DVDD:10667 0.02232
rDVDD/3592 DVDD:10663 DVDD:15710 0.0462825
rDVDD/3593 DVDD:10663 DVDD:10666 0.0603243
rDVDD/3594 DVDD:10663 DVDD:10664 0.5625
rDVDD/3595 DVDD:10659 DVDD:11177 0.02232
rDVDD/3596 DVDD:10659 DVDD:10753 0.02232
rDVDD/3597 DVDD:10658 DVDD:15763 0.0453096
rDVDD/3598 DVDD:10658 DVDD:10752 0.0589444
rDVDD/3599 DVDD:10658 DVDD:10659 0.5
rDVDD/3600 DVDD:9148 DVDD:13557 0.0117
rDVDD/3601 DVDD:9140 DVDD:13530 0.011682
rDVDD/3602 DVDD:9133 DVDD:9148 0.52
rDVDD/3603 DVDD:9132 DVDD:13242 0.01368
rDVDD/3604 DVDD:9132 DVDD:9133 0.433333
rDVDD/3605 DVDD:9125 DVDD:9140 0.52
rDVDD/3606 DVDD:9124 DVDD:13215 0.013662
rDVDD/3607 DVDD:9124 DVDD:9125 0.433333
rDVDD/3608 DVDD:9116 DVDD:9148 0.236776
rDVDD/3609 DVDD:9116 DVDD:9133 1.73333
rDVDD/3610 DVDD:9113 DVDD:9116 0.377206
rDVDD/3611 DVDD:9113 DVDD:9133 1.73333
rDVDD/3612 DVDD:9110 DVDD:9132 0.490893
rDVDD/3613 DVDD:9110 DVDD:9113 0.377206
rDVDD/3614 DVDD:9110 DVDD:9133 1.73333
rDVDD/3615 DVDD:9105 DVDD:9140 0.236794
rDVDD/3616 DVDD:9105 DVDD:9125 1.73333
rDVDD/3617 DVDD:9102 DVDD:9105 0.377206
rDVDD/3618 DVDD:9102 DVDD:9125 1.73333
rDVDD/3619 DVDD:9099 DVDD:9124 0.490911
rDVDD/3620 DVDD:9099 DVDD:9102 0.377206
rDVDD/3621 DVDD:9099 DVDD:9125 1.73333
rDVDD/3622 X52/X1/X2/X1/C0:pos DVDD:9125 3.65613
rDVDD/3623 X52/X1/X2/X1/C0:pos DVDD:9133 3.6566
rDVDD/3624 DVDD:9078 DVDD:9086 0.280062
rDVDD/3625 DVDD:9071 DVDD:9086 0.52
rDVDD/3626 DVDD:9070 DVDD:12927 0.01368
rDVDD/3627 DVDD:9070 DVDD:9071 0.433333
rDVDD/3628 DVDD:9063 DVDD:9078 0.52
rDVDD/3629 DVDD:9062 DVDD:12900 0.013662
rDVDD/3630 DVDD:9062 DVDD:9063 0.433333
rDVDD/3631 DVDD:9054 DVDD:9086 0.236776
rDVDD/3632 DVDD:9054 DVDD:9071 1.73333
rDVDD/3633 DVDD:9051 DVDD:9054 0.377206
rDVDD/3634 DVDD:9051 DVDD:9071 1.73333
rDVDD/3635 DVDD:9048 DVDD:9070 0.490893
rDVDD/3636 DVDD:9048 DVDD:9051 0.377206
rDVDD/3637 DVDD:9048 DVDD:9071 1.73333
rDVDD/3638 DVDD:9043 DVDD:9078 0.236794
rDVDD/3639 DVDD:9043 DVDD:9063 1.73333
rDVDD/3640 DVDD:9040 DVDD:9043 0.377206
rDVDD/3641 DVDD:9040 DVDD:9063 1.73333
rDVDD/3642 DVDD:9037 DVDD:9062 0.490911
rDVDD/3643 DVDD:9037 DVDD:9040 0.377206
rDVDD/3644 DVDD:9037 DVDD:9063 1.73333
rDVDD/3645 X52/X1/X2/X0/C0:pos DVDD:9063 3.65613
rDVDD/3646 X52/X1/X2/X0/C0:pos DVDD:9071 3.6566
rDVDD/3647 DVDD:8976 DVDD:12612 0.01368
rDVDD/3648 DVDD:8968 DVDD:12585 0.013662
rDVDD/3649 DVDD:8961 DVDD:8976 0.52
rDVDD/3650 DVDD:8960 DVDD:8961 0.433333
rDVDD/3651 DVDD:8953 DVDD:8968 0.52
rDVDD/3652 DVDD:8952 DVDD:8960 0.280062
rDVDD/3653 DVDD:8952 DVDD:8953 0.433333
rDVDD/3654 DVDD:8944 DVDD:8976 0.236776
rDVDD/3655 DVDD:8944 DVDD:8961 1.73333
rDVDD/3656 DVDD:8941 DVDD:8944 0.377206
rDVDD/3657 DVDD:8941 DVDD:8961 1.73333
rDVDD/3658 DVDD:8938 DVDD:8960 0.490893
rDVDD/3659 DVDD:8938 DVDD:8941 0.377206
rDVDD/3660 DVDD:8938 DVDD:8961 1.73333
rDVDD/3661 DVDD:8933 DVDD:8968 0.236794
rDVDD/3662 DVDD:8933 DVDD:8953 1.73333
rDVDD/3663 DVDD:8930 DVDD:8933 0.377206
rDVDD/3664 DVDD:8930 DVDD:8953 1.73333
rDVDD/3665 DVDD:8927 DVDD:8952 0.490911
rDVDD/3666 DVDD:8927 DVDD:8930 0.377206
rDVDD/3667 DVDD:8927 DVDD:8953 1.73333
rDVDD/3668 X52/X1/X1/X1/C0:pos DVDD:8953 3.65613
rDVDD/3669 X52/X1/X1/X1/C0:pos DVDD:8961 3.6566
rDVDD/3670 DVDD:8914 DVDD:12191 0.01368
rDVDD/3671 DVDD:8906 DVDD:12164 0.013662
rDVDD/3672 DVDD:8899 DVDD:8914 0.52
rDVDD/3673 DVDD:8898 DVDD:11527 0.00054
rDVDD/3674 DVDD:8898 DVDD:8899 0.433333
rDVDD/3675 DVDD:8891 DVDD:8906 0.52
rDVDD/3676 DVDD:8890 DVDD:11476 0.000522
rDVDD/3677 DVDD:8890 DVDD:8891 0.433333
rDVDD/3678 DVDD:8882 DVDD:8914 0.236776
rDVDD/3679 DVDD:8882 DVDD:8899 1.73333
rDVDD/3680 DVDD:8879 DVDD:8882 0.377206
rDVDD/3681 DVDD:8879 DVDD:8899 1.73333
rDVDD/3682 DVDD:8876 DVDD:8898 0.490893
rDVDD/3683 DVDD:8876 DVDD:8879 0.377206
rDVDD/3684 DVDD:8876 DVDD:8899 1.73333
rDVDD/3685 DVDD:8871 DVDD:8906 0.236794
rDVDD/3686 DVDD:8871 DVDD:8891 1.73333
rDVDD/3687 DVDD:8868 DVDD:8871 0.377206
rDVDD/3688 DVDD:8868 DVDD:8891 1.73333
rDVDD/3689 DVDD:8865 DVDD:8890 0.490911
rDVDD/3690 DVDD:8865 DVDD:8868 0.377206
rDVDD/3691 DVDD:8865 DVDD:8891 1.73333
rDVDD/3692 X52/X1/X1/X0/C0:pos DVDD:8891 3.65613
rDVDD/3693 X52/X1/X1/X0/C0:pos DVDD:8899 3.6566
rDVDD/3694 DVDD:8698 DVDD:13522 0.0117
rDVDD/3695 DVDD:8690 DVDD:13495 0.011682
rDVDD/3696 DVDD:8683 DVDD:8698 0.52
rDVDD/3697 DVDD:8682 DVDD:13207 0.01368
rDVDD/3698 DVDD:8682 DVDD:8683 0.433333
rDVDD/3699 DVDD:8675 DVDD:8690 0.52
rDVDD/3700 DVDD:8674 DVDD:13180 0.013662
rDVDD/3701 DVDD:8674 DVDD:8675 0.433333
rDVDD/3702 DVDD:8666 DVDD:8698 0.236776
rDVDD/3703 DVDD:8666 DVDD:8683 1.73333
rDVDD/3704 DVDD:8663 DVDD:8666 0.377206
rDVDD/3705 DVDD:8663 DVDD:8683 1.73333
rDVDD/3706 DVDD:8660 DVDD:8682 0.490893
rDVDD/3707 DVDD:8660 DVDD:8663 0.377206
rDVDD/3708 DVDD:8660 DVDD:8683 1.73333
rDVDD/3709 DVDD:8655 DVDD:8690 0.236794
rDVDD/3710 DVDD:8655 DVDD:8675 1.73333
rDVDD/3711 DVDD:8652 DVDD:8655 0.377206
rDVDD/3712 DVDD:8652 DVDD:8675 1.73333
rDVDD/3713 DVDD:8649 DVDD:8674 0.490911
rDVDD/3714 DVDD:8649 DVDD:8652 0.377206
rDVDD/3715 DVDD:8649 DVDD:8675 1.73333
rDVDD/3716 X52/X0/X2/X1/C0:pos DVDD:8675 3.65613
rDVDD/3717 X52/X0/X2/X1/C0:pos DVDD:8683 3.6566
rDVDD/3718 DVDD:8628 DVDD:8636 0.280062
rDVDD/3719 DVDD:8621 DVDD:8636 0.52
rDVDD/3720 DVDD:8620 DVDD:12892 0.01368
rDVDD/3721 DVDD:8620 DVDD:8621 0.433333
rDVDD/3722 DVDD:8613 DVDD:8628 0.52
rDVDD/3723 DVDD:8612 DVDD:12865 0.013662
rDVDD/3724 DVDD:8612 DVDD:8613 0.433333
rDVDD/3725 DVDD:8604 DVDD:8636 0.236776
rDVDD/3726 DVDD:8604 DVDD:8621 1.73333
rDVDD/3727 DVDD:8601 DVDD:8604 0.377206
rDVDD/3728 DVDD:8601 DVDD:8621 1.73333
rDVDD/3729 DVDD:8598 DVDD:8620 0.490893
rDVDD/3730 DVDD:8598 DVDD:8601 0.377206
rDVDD/3731 DVDD:8598 DVDD:8621 1.73333
rDVDD/3732 DVDD:8593 DVDD:8628 0.236794
rDVDD/3733 DVDD:8593 DVDD:8613 1.73333
rDVDD/3734 DVDD:8590 DVDD:8593 0.377206
rDVDD/3735 DVDD:8590 DVDD:8613 1.73333
rDVDD/3736 DVDD:8587 DVDD:8612 0.490911
rDVDD/3737 DVDD:8587 DVDD:8590 0.377206
rDVDD/3738 DVDD:8587 DVDD:8613 1.73333
rDVDD/3739 X52/X0/X2/X0/C0:pos DVDD:8613 3.65613
rDVDD/3740 X52/X0/X2/X0/C0:pos DVDD:8621 3.6566
rDVDD/3741 DVDD:8526 DVDD:12577 0.01368
rDVDD/3742 DVDD:8518 DVDD:12550 0.013662
rDVDD/3743 DVDD:8511 DVDD:8526 0.52
rDVDD/3744 DVDD:8510 DVDD:8511 0.433333
rDVDD/3745 DVDD:8503 DVDD:8518 0.52
rDVDD/3746 DVDD:8502 DVDD:8510 0.280062
rDVDD/3747 DVDD:8502 DVDD:8503 0.433333
rDVDD/3748 DVDD:8494 DVDD:8526 0.236776
rDVDD/3749 DVDD:8494 DVDD:8511 1.73333
rDVDD/3750 DVDD:8491 DVDD:8494 0.377206
rDVDD/3751 DVDD:8491 DVDD:8511 1.73333
rDVDD/3752 DVDD:8488 DVDD:8510 0.490893
rDVDD/3753 DVDD:8488 DVDD:8491 0.377206
rDVDD/3754 DVDD:8488 DVDD:8511 1.73333
rDVDD/3755 DVDD:8483 DVDD:8518 0.236794
rDVDD/3756 DVDD:8483 DVDD:8503 1.73333
rDVDD/3757 DVDD:8480 DVDD:8483 0.377206
rDVDD/3758 DVDD:8480 DVDD:8503 1.73333
rDVDD/3759 DVDD:8477 DVDD:8502 0.490911
rDVDD/3760 DVDD:8477 DVDD:8480 0.377206
rDVDD/3761 DVDD:8477 DVDD:8503 1.73333
rDVDD/3762 X52/X0/X1/X1/C0:pos DVDD:8503 3.65613
rDVDD/3763 X52/X0/X1/X1/C0:pos DVDD:8511 3.6566
rDVDD/3764 DVDD:8464 DVDD:12156 0.01368
rDVDD/3765 DVDD:8456 DVDD:12129 0.013662
rDVDD/3766 DVDD:8449 DVDD:8464 0.52
rDVDD/3767 DVDD:8448 DVDD:11468 0.00054
rDVDD/3768 DVDD:8448 DVDD:8449 0.433333
rDVDD/3769 DVDD:8441 DVDD:8456 0.52
rDVDD/3770 DVDD:8440 DVDD:11417 0.000522
rDVDD/3771 DVDD:8440 DVDD:8441 0.433333
rDVDD/3772 DVDD:8432 DVDD:8464 0.236776
rDVDD/3773 DVDD:8432 DVDD:8449 1.73333
rDVDD/3774 DVDD:8429 DVDD:8432 0.377206
rDVDD/3775 DVDD:8429 DVDD:8449 1.73333
rDVDD/3776 DVDD:8426 DVDD:8448 0.490893
rDVDD/3777 DVDD:8426 DVDD:8429 0.377206
rDVDD/3778 DVDD:8426 DVDD:8449 1.73333
rDVDD/3779 DVDD:8421 DVDD:8456 0.236794
rDVDD/3780 DVDD:8421 DVDD:8441 1.73333
rDVDD/3781 DVDD:8418 DVDD:8421 0.377206
rDVDD/3782 DVDD:8418 DVDD:8441 1.73333
rDVDD/3783 DVDD:8415 DVDD:8440 0.490911
rDVDD/3784 DVDD:8415 DVDD:8418 0.377206
rDVDD/3785 DVDD:8415 DVDD:8441 1.73333
rDVDD/3786 X52/X0/X1/X0/C0:pos DVDD:8441 3.65613
rDVDD/3787 X52/X0/X1/X0/C0:pos DVDD:8449 3.6566
rDVDD/3788 DVDD:8104 DVDD:13487 0.0117
rDVDD/3789 DVDD:8096 DVDD:13460 0.011682
rDVDD/3790 DVDD:8089 DVDD:8104 0.52
rDVDD/3791 DVDD:8088 DVDD:13172 0.01368
rDVDD/3792 DVDD:8088 DVDD:8089 0.433333
rDVDD/3793 DVDD:8081 DVDD:8096 0.52
rDVDD/3794 DVDD:8080 DVDD:13145 0.013662
rDVDD/3795 DVDD:8080 DVDD:8081 0.433333
rDVDD/3796 DVDD:8072 DVDD:8104 0.236776
rDVDD/3797 DVDD:8072 DVDD:8089 1.73333
rDVDD/3798 DVDD:8069 DVDD:8072 0.377206
rDVDD/3799 DVDD:8069 DVDD:8089 1.73333
rDVDD/3800 DVDD:8066 DVDD:8088 0.490893
rDVDD/3801 DVDD:8066 DVDD:8069 0.377206
rDVDD/3802 DVDD:8066 DVDD:8089 1.73333
rDVDD/3803 DVDD:8061 DVDD:8096 0.236794
rDVDD/3804 DVDD:8061 DVDD:8081 1.73333
rDVDD/3805 DVDD:8058 DVDD:8061 0.377206
rDVDD/3806 DVDD:8058 DVDD:8081 1.73333
rDVDD/3807 DVDD:8055 DVDD:8080 0.490911
rDVDD/3808 DVDD:8055 DVDD:8058 0.377206
rDVDD/3809 DVDD:8055 DVDD:8081 1.73333
rDVDD/3810 X51/X1/X2/X1/C0:pos DVDD:8081 3.65613
rDVDD/3811 X51/X1/X2/X1/C0:pos DVDD:8089 3.6566
rDVDD/3812 DVDD:8034 DVDD:8042 0.280062
rDVDD/3813 DVDD:8027 DVDD:8042 0.52
rDVDD/3814 DVDD:8026 DVDD:12857 0.01368
rDVDD/3815 DVDD:8026 DVDD:8027 0.433333
rDVDD/3816 DVDD:8019 DVDD:8034 0.52
rDVDD/3817 DVDD:8018 DVDD:12830 0.013662
rDVDD/3818 DVDD:8018 DVDD:8019 0.433333
rDVDD/3819 DVDD:8010 DVDD:8042 0.236776
rDVDD/3820 DVDD:8010 DVDD:8027 1.73333
rDVDD/3821 DVDD:8007 DVDD:8010 0.377206
rDVDD/3822 DVDD:8007 DVDD:8027 1.73333
rDVDD/3823 DVDD:8004 DVDD:8026 0.490893
rDVDD/3824 DVDD:8004 DVDD:8007 0.377206
rDVDD/3825 DVDD:8004 DVDD:8027 1.73333
rDVDD/3826 DVDD:7999 DVDD:8034 0.236794
rDVDD/3827 DVDD:7999 DVDD:8019 1.73333
rDVDD/3828 DVDD:7996 DVDD:7999 0.377206
rDVDD/3829 DVDD:7996 DVDD:8019 1.73333
rDVDD/3830 DVDD:7993 DVDD:8018 0.490911
rDVDD/3831 DVDD:7993 DVDD:7996 0.377206
rDVDD/3832 DVDD:7993 DVDD:8019 1.73333
rDVDD/3833 X51/X1/X2/X0/C0:pos DVDD:8019 3.65613
rDVDD/3834 X51/X1/X2/X0/C0:pos DVDD:8027 3.6566
rDVDD/3835 DVDD:7932 DVDD:12542 0.01368
rDVDD/3836 DVDD:7924 DVDD:12515 0.013662
rDVDD/3837 DVDD:7917 DVDD:7932 0.52
rDVDD/3838 DVDD:7916 DVDD:7917 0.433333
rDVDD/3839 DVDD:7909 DVDD:7924 0.52
rDVDD/3840 DVDD:7908 DVDD:7916 0.280062
rDVDD/3841 DVDD:7908 DVDD:7909 0.433333
rDVDD/3842 DVDD:7900 DVDD:7932 0.236776
rDVDD/3843 DVDD:7900 DVDD:7917 1.73333
rDVDD/3844 DVDD:7897 DVDD:7900 0.377206
rDVDD/3845 DVDD:7897 DVDD:7917 1.73333
rDVDD/3846 DVDD:7894 DVDD:7916 0.490893
rDVDD/3847 DVDD:7894 DVDD:7897 0.377206
rDVDD/3848 DVDD:7894 DVDD:7917 1.73333
rDVDD/3849 DVDD:7889 DVDD:7924 0.236794
rDVDD/3850 DVDD:7889 DVDD:7909 1.73333
rDVDD/3851 DVDD:7886 DVDD:7889 0.377206
rDVDD/3852 DVDD:7886 DVDD:7909 1.73333
rDVDD/3853 DVDD:7883 DVDD:7908 0.490911
rDVDD/3854 DVDD:7883 DVDD:7886 0.377206
rDVDD/3855 DVDD:7883 DVDD:7909 1.73333
rDVDD/3856 X51/X1/X1/X1/C0:pos DVDD:7909 3.65613
rDVDD/3857 X51/X1/X1/X1/C0:pos DVDD:7917 3.6566
rDVDD/3858 DVDD:7870 DVDD:12121 0.01368
rDVDD/3859 DVDD:7862 DVDD:12094 0.013662
rDVDD/3860 DVDD:7855 DVDD:7870 0.52
rDVDD/3861 DVDD:7854 DVDD:11409 0.00054
rDVDD/3862 DVDD:7854 DVDD:7855 0.433333
rDVDD/3863 DVDD:7847 DVDD:7862 0.52
rDVDD/3864 DVDD:7846 DVDD:11358 0.000522
rDVDD/3865 DVDD:7846 DVDD:7847 0.433333
rDVDD/3866 DVDD:7838 DVDD:7870 0.236776
rDVDD/3867 DVDD:7838 DVDD:7855 1.73333
rDVDD/3868 DVDD:7835 DVDD:7838 0.377206
rDVDD/3869 DVDD:7835 DVDD:7855 1.73333
rDVDD/3870 DVDD:7832 DVDD:7854 0.490893
rDVDD/3871 DVDD:7832 DVDD:7835 0.377206
rDVDD/3872 DVDD:7832 DVDD:7855 1.73333
rDVDD/3873 DVDD:7827 DVDD:7862 0.236794
rDVDD/3874 DVDD:7827 DVDD:7847 1.73333
rDVDD/3875 DVDD:7824 DVDD:7827 0.377206
rDVDD/3876 DVDD:7824 DVDD:7847 1.73333
rDVDD/3877 DVDD:7821 DVDD:7846 0.490911
rDVDD/3878 DVDD:7821 DVDD:7824 0.377206
rDVDD/3879 DVDD:7821 DVDD:7847 1.73333
rDVDD/3880 X51/X1/X1/X0/C0:pos DVDD:7847 3.65613
rDVDD/3881 X51/X1/X1/X0/C0:pos DVDD:7855 3.6566
rDVDD/3882 DVDD:7654 DVDD:13452 0.0117
rDVDD/3883 DVDD:7646 DVDD:13425 0.011682
rDVDD/3884 DVDD:7639 DVDD:7654 0.52
rDVDD/3885 DVDD:7638 DVDD:13137 0.01368
rDVDD/3886 DVDD:7638 DVDD:7639 0.433333
rDVDD/3887 DVDD:7631 DVDD:7646 0.52
rDVDD/3888 DVDD:7630 DVDD:13110 0.013662
rDVDD/3889 DVDD:7630 DVDD:7631 0.433333
rDVDD/3890 DVDD:7622 DVDD:7654 0.236776
rDVDD/3891 DVDD:7622 DVDD:7639 1.73333
rDVDD/3892 DVDD:7619 DVDD:7622 0.377206
rDVDD/3893 DVDD:7619 DVDD:7639 1.73333
rDVDD/3894 DVDD:7616 DVDD:7638 0.490893
rDVDD/3895 DVDD:7616 DVDD:7619 0.377206
rDVDD/3896 DVDD:7616 DVDD:7639 1.73333
rDVDD/3897 DVDD:7611 DVDD:7646 0.236794
rDVDD/3898 DVDD:7611 DVDD:7631 1.73333
rDVDD/3899 DVDD:7608 DVDD:7611 0.377206
rDVDD/3900 DVDD:7608 DVDD:7631 1.73333
rDVDD/3901 DVDD:7605 DVDD:7630 0.490911
rDVDD/3902 DVDD:7605 DVDD:7608 0.377206
rDVDD/3903 DVDD:7605 DVDD:7631 1.73333
rDVDD/3904 X51/X0/X2/X1/C0:pos DVDD:7631 3.65613
rDVDD/3905 X51/X0/X2/X1/C0:pos DVDD:7639 3.6566
rDVDD/3906 DVDD:7584 DVDD:7592 0.280062
rDVDD/3907 DVDD:7577 DVDD:7592 0.52
rDVDD/3908 DVDD:7576 DVDD:12822 0.01368
rDVDD/3909 DVDD:7576 DVDD:7577 0.433333
rDVDD/3910 DVDD:7569 DVDD:7584 0.52
rDVDD/3911 DVDD:7568 DVDD:12795 0.013662
rDVDD/3912 DVDD:7568 DVDD:7569 0.433333
rDVDD/3913 DVDD:7560 DVDD:7592 0.236776
rDVDD/3914 DVDD:7560 DVDD:7577 1.73333
rDVDD/3915 DVDD:7557 DVDD:7560 0.377206
rDVDD/3916 DVDD:7557 DVDD:7577 1.73333
rDVDD/3917 DVDD:7554 DVDD:7576 0.490893
rDVDD/3918 DVDD:7554 DVDD:7557 0.377206
rDVDD/3919 DVDD:7554 DVDD:7577 1.73333
rDVDD/3920 DVDD:7549 DVDD:7584 0.236794
rDVDD/3921 DVDD:7549 DVDD:7569 1.73333
rDVDD/3922 DVDD:7546 DVDD:7549 0.377206
rDVDD/3923 DVDD:7546 DVDD:7569 1.73333
rDVDD/3924 DVDD:7543 DVDD:7568 0.490911
rDVDD/3925 DVDD:7543 DVDD:7546 0.377206
rDVDD/3926 DVDD:7543 DVDD:7569 1.73333
rDVDD/3927 X51/X0/X2/X0/C0:pos DVDD:7569 3.65613
rDVDD/3928 X51/X0/X2/X0/C0:pos DVDD:7577 3.6566
rDVDD/3929 DVDD:7482 DVDD:12507 0.01368
rDVDD/3930 DVDD:7474 DVDD:12480 0.013662
rDVDD/3931 DVDD:7467 DVDD:7482 0.52
rDVDD/3932 DVDD:7466 DVDD:7467 0.433333
rDVDD/3933 DVDD:7459 DVDD:7474 0.52
rDVDD/3934 DVDD:7458 DVDD:7466 0.280062
rDVDD/3935 DVDD:7458 DVDD:7459 0.433333
rDVDD/3936 DVDD:7450 DVDD:7482 0.236776
rDVDD/3937 DVDD:7450 DVDD:7467 1.73333
rDVDD/3938 DVDD:7447 DVDD:7450 0.377206
rDVDD/3939 DVDD:7447 DVDD:7467 1.73333
rDVDD/3940 DVDD:7444 DVDD:7466 0.490893
rDVDD/3941 DVDD:7444 DVDD:7447 0.377206
rDVDD/3942 DVDD:7444 DVDD:7467 1.73333
rDVDD/3943 DVDD:7439 DVDD:7474 0.236794
rDVDD/3944 DVDD:7439 DVDD:7459 1.73333
rDVDD/3945 DVDD:7436 DVDD:7439 0.377206
rDVDD/3946 DVDD:7436 DVDD:7459 1.73333
rDVDD/3947 DVDD:7433 DVDD:7458 0.490911
rDVDD/3948 DVDD:7433 DVDD:7436 0.377206
rDVDD/3949 DVDD:7433 DVDD:7459 1.73333
rDVDD/3950 X51/X0/X1/X1/C0:pos DVDD:7459 3.65613
rDVDD/3951 X51/X0/X1/X1/C0:pos DVDD:7467 3.6566
rDVDD/3952 DVDD:7420 DVDD:12086 0.01368
rDVDD/3953 DVDD:7412 DVDD:12059 0.013662
rDVDD/3954 DVDD:7405 DVDD:7420 0.52
rDVDD/3955 DVDD:7404 DVDD:11350 0.00054
rDVDD/3956 DVDD:7404 DVDD:7405 0.433333
rDVDD/3957 DVDD:7397 DVDD:7412 0.52
rDVDD/3958 DVDD:7396 DVDD:11299 0.000522
rDVDD/3959 DVDD:7396 DVDD:7397 0.433333
rDVDD/3960 DVDD:7388 DVDD:7420 0.236776
rDVDD/3961 DVDD:7388 DVDD:7405 1.73333
rDVDD/3962 DVDD:7385 DVDD:7388 0.377206
rDVDD/3963 DVDD:7385 DVDD:7405 1.73333
rDVDD/3964 DVDD:7382 DVDD:7404 0.490893
rDVDD/3965 DVDD:7382 DVDD:7385 0.377206
rDVDD/3966 DVDD:7382 DVDD:7405 1.73333
rDVDD/3967 DVDD:7377 DVDD:7412 0.236794
rDVDD/3968 DVDD:7377 DVDD:7397 1.73333
rDVDD/3969 DVDD:7374 DVDD:7377 0.377206
rDVDD/3970 DVDD:7374 DVDD:7397 1.73333
rDVDD/3971 DVDD:7371 DVDD:7396 0.490911
rDVDD/3972 DVDD:7371 DVDD:7374 0.377206
rDVDD/3973 DVDD:7371 DVDD:7397 1.73333
rDVDD/3974 X51/X0/X1/X0/C0:pos DVDD:7397 3.65613
rDVDD/3975 X51/X0/X1/X0/C0:pos DVDD:7405 3.6566
rDVDD/3976 DVDD:7060 DVDD:13417 0.0117
rDVDD/3977 DVDD:7052 DVDD:13390 0.011682
rDVDD/3978 DVDD:7045 DVDD:7060 0.52
rDVDD/3979 DVDD:7044 DVDD:13102 0.01368
rDVDD/3980 DVDD:7044 DVDD:7045 0.433333
rDVDD/3981 DVDD:7037 DVDD:7052 0.52
rDVDD/3982 DVDD:7036 DVDD:13075 0.013662
rDVDD/3983 DVDD:7036 DVDD:7037 0.433333
rDVDD/3984 DVDD:7028 DVDD:7060 0.236776
rDVDD/3985 DVDD:7028 DVDD:7045 1.73333
rDVDD/3986 DVDD:7025 DVDD:7028 0.377206
rDVDD/3987 DVDD:7025 DVDD:7045 1.73333
rDVDD/3988 DVDD:7022 DVDD:7044 0.490893
rDVDD/3989 DVDD:7022 DVDD:7025 0.377206
rDVDD/3990 DVDD:7022 DVDD:7045 1.73333
rDVDD/3991 DVDD:7017 DVDD:7052 0.236794
rDVDD/3992 DVDD:7017 DVDD:7037 1.73333
rDVDD/3993 DVDD:7014 DVDD:7017 0.377206
rDVDD/3994 DVDD:7014 DVDD:7037 1.73333
rDVDD/3995 DVDD:7011 DVDD:7036 0.490911
rDVDD/3996 DVDD:7011 DVDD:7014 0.377206
rDVDD/3997 DVDD:7011 DVDD:7037 1.73333
rDVDD/3998 X50/X1/X2/X1/C0:pos DVDD:7037 3.65613
rDVDD/3999 X50/X1/X2/X1/C0:pos DVDD:7045 3.6566
rDVDD/4000 DVDD:6990 DVDD:6998 0.280062
rDVDD/4001 DVDD:6983 DVDD:6998 0.52
rDVDD/4002 DVDD:6982 DVDD:12787 0.01368
rDVDD/4003 DVDD:6982 DVDD:6983 0.433333
rDVDD/4004 DVDD:6975 DVDD:6990 0.52
rDVDD/4005 DVDD:6974 DVDD:12760 0.013662
rDVDD/4006 DVDD:6974 DVDD:6975 0.433333
rDVDD/4007 DVDD:6966 DVDD:6998 0.236776
rDVDD/4008 DVDD:6966 DVDD:6983 1.73333
rDVDD/4009 DVDD:6963 DVDD:6966 0.377206
rDVDD/4010 DVDD:6963 DVDD:6983 1.73333
rDVDD/4011 DVDD:6960 DVDD:6982 0.490893
rDVDD/4012 DVDD:6960 DVDD:6963 0.377206
rDVDD/4013 DVDD:6960 DVDD:6983 1.73333
rDVDD/4014 DVDD:6955 DVDD:6990 0.236794
rDVDD/4015 DVDD:6955 DVDD:6975 1.73333
rDVDD/4016 DVDD:6952 DVDD:6955 0.377206
rDVDD/4017 DVDD:6952 DVDD:6975 1.73333
rDVDD/4018 DVDD:6949 DVDD:6974 0.490911
rDVDD/4019 DVDD:6949 DVDD:6952 0.377206
rDVDD/4020 DVDD:6949 DVDD:6975 1.73333
rDVDD/4021 X50/X1/X2/X0/C0:pos DVDD:6975 3.65613
rDVDD/4022 X50/X1/X2/X0/C0:pos DVDD:6983 3.6566
rDVDD/4023 DVDD:6888 DVDD:12472 0.01368
rDVDD/4024 DVDD:6880 DVDD:12445 0.013662
rDVDD/4025 DVDD:6873 DVDD:6888 0.52
rDVDD/4026 DVDD:6872 DVDD:6873 0.433333
rDVDD/4027 DVDD:6865 DVDD:6880 0.52
rDVDD/4028 DVDD:6864 DVDD:6872 0.280062
rDVDD/4029 DVDD:6864 DVDD:6865 0.433333
rDVDD/4030 DVDD:6856 DVDD:6888 0.236776
rDVDD/4031 DVDD:6856 DVDD:6873 1.73333
rDVDD/4032 DVDD:6853 DVDD:6856 0.377206
rDVDD/4033 DVDD:6853 DVDD:6873 1.73333
rDVDD/4034 DVDD:6850 DVDD:6872 0.490893
rDVDD/4035 DVDD:6850 DVDD:6853 0.377206
rDVDD/4036 DVDD:6850 DVDD:6873 1.73333
rDVDD/4037 DVDD:6845 DVDD:6880 0.236794
rDVDD/4038 DVDD:6845 DVDD:6865 1.73333
rDVDD/4039 DVDD:6842 DVDD:6845 0.377206
rDVDD/4040 DVDD:6842 DVDD:6865 1.73333
rDVDD/4041 DVDD:6839 DVDD:6864 0.490911
rDVDD/4042 DVDD:6839 DVDD:6842 0.377206
rDVDD/4043 DVDD:6839 DVDD:6865 1.73333
rDVDD/4044 X50/X1/X1/X1/C0:pos DVDD:6865 3.65613
rDVDD/4045 X50/X1/X1/X1/C0:pos DVDD:6873 3.6566
rDVDD/4046 DVDD:6826 DVDD:12051 0.01368
rDVDD/4047 DVDD:6818 DVDD:12024 0.013662
rDVDD/4048 DVDD:6811 DVDD:6826 0.52
rDVDD/4049 DVDD:6810 DVDD:10767 0.00054
rDVDD/4050 DVDD:6810 DVDD:6811 0.433333
rDVDD/4051 DVDD:6803 DVDD:6818 0.52
rDVDD/4052 DVDD:6802 DVDD:10762 0.000522
rDVDD/4053 DVDD:6802 DVDD:6803 0.433333
rDVDD/4054 DVDD:6794 DVDD:6826 0.236776
rDVDD/4055 DVDD:6794 DVDD:6811 1.73333
rDVDD/4056 DVDD:6791 DVDD:6794 0.377206
rDVDD/4057 DVDD:6791 DVDD:6811 1.73333
rDVDD/4058 DVDD:6788 DVDD:6810 0.490893
rDVDD/4059 DVDD:6788 DVDD:6791 0.377206
rDVDD/4060 DVDD:6788 DVDD:6811 1.73333
rDVDD/4061 DVDD:6783 DVDD:6818 0.236794
rDVDD/4062 DVDD:6783 DVDD:6803 1.73333
rDVDD/4063 DVDD:6780 DVDD:6783 0.377206
rDVDD/4064 DVDD:6780 DVDD:6803 1.73333
rDVDD/4065 DVDD:6777 DVDD:6802 0.490911
rDVDD/4066 DVDD:6777 DVDD:6780 0.377206
rDVDD/4067 DVDD:6777 DVDD:6803 1.73333
rDVDD/4068 X50/X1/X1/X0/C0:pos DVDD:6803 3.65613
rDVDD/4069 X50/X1/X1/X0/C0:pos DVDD:6811 3.6566
rDVDD/4070 DVDD:6610 DVDD:13382 0.0117
rDVDD/4071 DVDD:6602 DVDD:13355 0.011682
rDVDD/4072 DVDD:6595 DVDD:6610 0.52
rDVDD/4073 DVDD:6594 DVDD:13067 0.01368
rDVDD/4074 DVDD:6594 DVDD:6595 0.433333
rDVDD/4075 DVDD:6587 DVDD:6602 0.52
rDVDD/4076 DVDD:6586 DVDD:13040 0.013662
rDVDD/4077 DVDD:6586 DVDD:6587 0.433333
rDVDD/4078 DVDD:6578 DVDD:6610 0.236776
rDVDD/4079 DVDD:6578 DVDD:6595 1.73333
rDVDD/4080 DVDD:6575 DVDD:6578 0.377206
rDVDD/4081 DVDD:6575 DVDD:6595 1.73333
rDVDD/4082 DVDD:6572 DVDD:6594 0.490893
rDVDD/4083 DVDD:6572 DVDD:6575 0.377206
rDVDD/4084 DVDD:6572 DVDD:6595 1.73333
rDVDD/4085 DVDD:6567 DVDD:6602 0.236794
rDVDD/4086 DVDD:6567 DVDD:6587 1.73333
rDVDD/4087 DVDD:6564 DVDD:6567 0.377206
rDVDD/4088 DVDD:6564 DVDD:6587 1.73333
rDVDD/4089 DVDD:6561 DVDD:6586 0.490911
rDVDD/4090 DVDD:6561 DVDD:6564 0.377206
rDVDD/4091 DVDD:6561 DVDD:6587 1.73333
rDVDD/4092 X50/X0/X2/X1/C0:pos DVDD:6587 3.65613
rDVDD/4093 X50/X0/X2/X1/C0:pos DVDD:6595 3.6566
rDVDD/4094 DVDD:6540 DVDD:6548 0.280062
rDVDD/4095 DVDD:6533 DVDD:6548 0.52
rDVDD/4096 DVDD:6532 DVDD:12752 0.01368
rDVDD/4097 DVDD:6532 DVDD:6533 0.433333
rDVDD/4098 DVDD:6525 DVDD:6540 0.52
rDVDD/4099 DVDD:6524 DVDD:12725 0.013662
rDVDD/4100 DVDD:6524 DVDD:6525 0.433333
rDVDD/4101 DVDD:6516 DVDD:6548 0.236776
rDVDD/4102 DVDD:6516 DVDD:6533 1.73333
rDVDD/4103 DVDD:6513 DVDD:6516 0.377206
rDVDD/4104 DVDD:6513 DVDD:6533 1.73333
rDVDD/4105 DVDD:6510 DVDD:6532 0.490893
rDVDD/4106 DVDD:6510 DVDD:6513 0.377206
rDVDD/4107 DVDD:6510 DVDD:6533 1.73333
rDVDD/4108 DVDD:6505 DVDD:6540 0.236794
rDVDD/4109 DVDD:6505 DVDD:6525 1.73333
rDVDD/4110 DVDD:6502 DVDD:6505 0.377206
rDVDD/4111 DVDD:6502 DVDD:6525 1.73333
rDVDD/4112 DVDD:6499 DVDD:6524 0.490911
rDVDD/4113 DVDD:6499 DVDD:6502 0.377206
rDVDD/4114 DVDD:6499 DVDD:6525 1.73333
rDVDD/4115 X50/X0/X2/X0/C0:pos DVDD:6525 3.65613
rDVDD/4116 X50/X0/X2/X0/C0:pos DVDD:6533 3.6566
rDVDD/4117 DVDD:6438 DVDD:12437 0.01368
rDVDD/4118 DVDD:6430 DVDD:12410 0.013662
rDVDD/4119 DVDD:6423 DVDD:6438 0.52
rDVDD/4120 DVDD:6422 DVDD:6423 0.433333
rDVDD/4121 DVDD:6415 DVDD:6430 0.52
rDVDD/4122 DVDD:6414 DVDD:6422 0.280062
rDVDD/4123 DVDD:6414 DVDD:6415 0.433333
rDVDD/4124 DVDD:6406 DVDD:6438 0.236776
rDVDD/4125 DVDD:6406 DVDD:6423 1.73333
rDVDD/4126 DVDD:6403 DVDD:6406 0.377206
rDVDD/4127 DVDD:6403 DVDD:6423 1.73333
rDVDD/4128 DVDD:6400 DVDD:6422 0.490893
rDVDD/4129 DVDD:6400 DVDD:6403 0.377206
rDVDD/4130 DVDD:6400 DVDD:6423 1.73333
rDVDD/4131 DVDD:6395 DVDD:6430 0.236794
rDVDD/4132 DVDD:6395 DVDD:6415 1.73333
rDVDD/4133 DVDD:6392 DVDD:6395 0.377206
rDVDD/4134 DVDD:6392 DVDD:6415 1.73333
rDVDD/4135 DVDD:6389 DVDD:6414 0.490911
rDVDD/4136 DVDD:6389 DVDD:6392 0.377206
rDVDD/4137 DVDD:6389 DVDD:6415 1.73333
rDVDD/4138 X50/X0/X1/X1/C0:pos DVDD:6415 3.65613
rDVDD/4139 X50/X0/X1/X1/C0:pos DVDD:6423 3.6566
rDVDD/4140 DVDD:6376 DVDD:12016 0.01368
rDVDD/4141 DVDD:6368 DVDD:11989 0.013662
rDVDD/4142 DVDD:6361 DVDD:6376 0.52
rDVDD/4143 DVDD:6360 DVDD:11248 0.00054
rDVDD/4144 DVDD:6360 DVDD:6361 0.433333
rDVDD/4145 DVDD:6353 DVDD:6368 0.52
rDVDD/4146 DVDD:6352 DVDD:11222 0.011682
rDVDD/4147 DVDD:6352 DVDD:6353 0.433333
rDVDD/4148 DVDD:6344 DVDD:6376 0.236776
rDVDD/4149 DVDD:6344 DVDD:6361 1.73333
rDVDD/4150 DVDD:6341 DVDD:6344 0.377206
rDVDD/4151 DVDD:6341 DVDD:6361 1.73333
rDVDD/4152 DVDD:6338 DVDD:6360 0.490893
rDVDD/4153 DVDD:6338 DVDD:6341 0.377206
rDVDD/4154 DVDD:6338 DVDD:6361 1.73333
rDVDD/4155 DVDD:6333 DVDD:6368 0.236794
rDVDD/4156 DVDD:6333 DVDD:6353 1.73333
rDVDD/4157 DVDD:6330 DVDD:6333 0.377206
rDVDD/4158 DVDD:6330 DVDD:6353 1.73333
rDVDD/4159 DVDD:6327 DVDD:6352 0.490911
rDVDD/4160 DVDD:6327 DVDD:6330 0.377206
rDVDD/4161 DVDD:6327 DVDD:6353 1.73333
rDVDD/4162 X50/X0/X1/X0/C0:pos DVDD:6353 3.65613
rDVDD/4163 X50/X0/X1/X0/C0:pos DVDD:6361 3.6566
rDVDD/4164 DVDD:6016 DVDD:13347 0.0117
rDVDD/4165 DVDD:6008 DVDD:13320 0.011682
rDVDD/4166 DVDD:6001 DVDD:6016 0.52
rDVDD/4167 DVDD:6000 DVDD:13032 0.01368
rDVDD/4168 DVDD:6000 DVDD:6001 0.433333
rDVDD/4169 DVDD:5993 DVDD:6008 0.52
rDVDD/4170 DVDD:5992 DVDD:13005 0.013662
rDVDD/4171 DVDD:5992 DVDD:5993 0.433333
rDVDD/4172 DVDD:5984 DVDD:6016 0.236776
rDVDD/4173 DVDD:5984 DVDD:6001 1.73333
rDVDD/4174 DVDD:5981 DVDD:5984 0.377206
rDVDD/4175 DVDD:5981 DVDD:6001 1.73333
rDVDD/4176 DVDD:5978 DVDD:6000 0.490893
rDVDD/4177 DVDD:5978 DVDD:5981 0.377206
rDVDD/4178 DVDD:5978 DVDD:6001 1.73333
rDVDD/4179 DVDD:5973 DVDD:6008 0.236794
rDVDD/4180 DVDD:5973 DVDD:5993 1.73333
rDVDD/4181 DVDD:5970 DVDD:5973 0.377206
rDVDD/4182 DVDD:5970 DVDD:5993 1.73333
rDVDD/4183 DVDD:5967 DVDD:5992 0.490911
rDVDD/4184 DVDD:5967 DVDD:5970 0.377206
rDVDD/4185 DVDD:5967 DVDD:5993 1.73333
rDVDD/4186 X49/X1/X2/X1/C0:pos DVDD:5993 3.65613
rDVDD/4187 X49/X1/X2/X1/C0:pos DVDD:6001 3.6566
rDVDD/4188 DVDD:5946 DVDD:5954 0.280062
rDVDD/4189 DVDD:5939 DVDD:5954 0.52
rDVDD/4190 DVDD:5938 DVDD:12717 0.01368
rDVDD/4191 DVDD:5938 DVDD:5939 0.433333
rDVDD/4192 DVDD:5931 DVDD:5946 0.52
rDVDD/4193 DVDD:5930 DVDD:12690 0.013662
rDVDD/4194 DVDD:5930 DVDD:5931 0.433333
rDVDD/4195 DVDD:5922 DVDD:5954 0.236776
rDVDD/4196 DVDD:5922 DVDD:5939 1.73333
rDVDD/4197 DVDD:5919 DVDD:5922 0.377206
rDVDD/4198 DVDD:5919 DVDD:5939 1.73333
rDVDD/4199 DVDD:5916 DVDD:5938 0.490893
rDVDD/4200 DVDD:5916 DVDD:5919 0.377206
rDVDD/4201 DVDD:5916 DVDD:5939 1.73333
rDVDD/4202 DVDD:5911 DVDD:5946 0.236794
rDVDD/4203 DVDD:5911 DVDD:5931 1.73333
rDVDD/4204 DVDD:5908 DVDD:5911 0.377206
rDVDD/4205 DVDD:5908 DVDD:5931 1.73333
rDVDD/4206 DVDD:5905 DVDD:5930 0.490911
rDVDD/4207 DVDD:5905 DVDD:5908 0.377206
rDVDD/4208 DVDD:5905 DVDD:5931 1.73333
rDVDD/4209 X49/X1/X2/X0/C0:pos DVDD:5931 3.65613
rDVDD/4210 X49/X1/X2/X0/C0:pos DVDD:5939 3.6566
rDVDD/4211 DVDD:5844 DVDD:12402 0.01368
rDVDD/4212 DVDD:5836 DVDD:12375 0.013662
rDVDD/4213 DVDD:5829 DVDD:5844 0.52
rDVDD/4214 DVDD:5828 DVDD:5829 0.433333
rDVDD/4215 DVDD:5821 DVDD:5836 0.52
rDVDD/4216 DVDD:5820 DVDD:5828 0.280062
rDVDD/4217 DVDD:5820 DVDD:5821 0.433333
rDVDD/4218 DVDD:5812 DVDD:5844 0.236776
rDVDD/4219 DVDD:5812 DVDD:5829 1.73333
rDVDD/4220 DVDD:5809 DVDD:5812 0.377206
rDVDD/4221 DVDD:5809 DVDD:5829 1.73333
rDVDD/4222 DVDD:5806 DVDD:5828 0.490893
rDVDD/4223 DVDD:5806 DVDD:5809 0.377206
rDVDD/4224 DVDD:5806 DVDD:5829 1.73333
rDVDD/4225 DVDD:5801 DVDD:5836 0.236794
rDVDD/4226 DVDD:5801 DVDD:5821 1.73333
rDVDD/4227 DVDD:5798 DVDD:5801 0.377206
rDVDD/4228 DVDD:5798 DVDD:5821 1.73333
rDVDD/4229 DVDD:5795 DVDD:5820 0.490911
rDVDD/4230 DVDD:5795 DVDD:5798 0.377206
rDVDD/4231 DVDD:5795 DVDD:5821 1.73333
rDVDD/4232 X49/X1/X1/X1/C0:pos DVDD:5821 3.65613
rDVDD/4233 X49/X1/X1/X1/C0:pos DVDD:5829 3.6566
rDVDD/4234 DVDD:5782 DVDD:11981 0.01368
rDVDD/4235 DVDD:5774 DVDD:11954 0.013662
rDVDD/4236 DVDD:5767 DVDD:5782 0.52
rDVDD/4237 DVDD:5766 DVDD:11214 0.00054
rDVDD/4238 DVDD:5766 DVDD:5767 0.433333
rDVDD/4239 DVDD:5759 DVDD:5774 0.52
rDVDD/4240 DVDD:5758 DVDD:11196 0.011682
rDVDD/4241 DVDD:5758 DVDD:5759 0.433333
rDVDD/4242 DVDD:5750 DVDD:5782 0.236776
rDVDD/4243 DVDD:5750 DVDD:5767 1.73333
rDVDD/4244 DVDD:5747 DVDD:5750 0.377206
rDVDD/4245 DVDD:5747 DVDD:5767 1.73333
rDVDD/4246 DVDD:5744 DVDD:5766 0.490893
rDVDD/4247 DVDD:5744 DVDD:5747 0.377206
rDVDD/4248 DVDD:5744 DVDD:5767 1.73333
rDVDD/4249 DVDD:5739 DVDD:5774 0.236794
rDVDD/4250 DVDD:5739 DVDD:5759 1.73333
rDVDD/4251 DVDD:5736 DVDD:5739 0.377206
rDVDD/4252 DVDD:5736 DVDD:5759 1.73333
rDVDD/4253 DVDD:5733 DVDD:5758 0.490911
rDVDD/4254 DVDD:5733 DVDD:5736 0.377206
rDVDD/4255 DVDD:5733 DVDD:5759 1.73333
rDVDD/4256 X49/X1/X1/X0/C0:pos DVDD:5759 3.65613
rDVDD/4257 X49/X1/X1/X0/C0:pos DVDD:5767 3.6566
rDVDD/4258 DVDD:5566 DVDD:13312 0.0117
rDVDD/4259 DVDD:5558 DVDD:13285 0.011682
rDVDD/4260 DVDD:5551 DVDD:5566 0.52
rDVDD/4261 DVDD:5550 DVDD:12997 0.01368
rDVDD/4262 DVDD:5550 DVDD:5551 0.433333
rDVDD/4263 DVDD:5543 DVDD:5558 0.52
rDVDD/4264 DVDD:5542 DVDD:12970 0.013662
rDVDD/4265 DVDD:5542 DVDD:5543 0.433333
rDVDD/4266 DVDD:5534 DVDD:5566 0.236776
rDVDD/4267 DVDD:5534 DVDD:5551 1.73333
rDVDD/4268 DVDD:5531 DVDD:5534 0.377206
rDVDD/4269 DVDD:5531 DVDD:5551 1.73333
rDVDD/4270 DVDD:5528 DVDD:5550 0.490893
rDVDD/4271 DVDD:5528 DVDD:5531 0.377206
rDVDD/4272 DVDD:5528 DVDD:5551 1.73333
rDVDD/4273 DVDD:5523 DVDD:5558 0.236794
rDVDD/4274 DVDD:5523 DVDD:5543 1.73333
rDVDD/4275 DVDD:5520 DVDD:5523 0.377206
rDVDD/4276 DVDD:5520 DVDD:5543 1.73333
rDVDD/4277 DVDD:5517 DVDD:5542 0.490911
rDVDD/4278 DVDD:5517 DVDD:5520 0.377206
rDVDD/4279 DVDD:5517 DVDD:5543 1.73333
rDVDD/4280 X49/X0/X2/X1/C0:pos DVDD:5543 3.65613
rDVDD/4281 X49/X0/X2/X1/C0:pos DVDD:5551 3.6566
rDVDD/4282 DVDD:5496 DVDD:5504 0.280062
rDVDD/4283 DVDD:5489 DVDD:5504 0.52
rDVDD/4284 DVDD:5488 DVDD:12682 0.01368
rDVDD/4285 DVDD:5488 DVDD:5489 0.433333
rDVDD/4286 DVDD:5481 DVDD:5496 0.52
rDVDD/4287 DVDD:5480 DVDD:12655 0.013662
rDVDD/4288 DVDD:5480 DVDD:5481 0.433333
rDVDD/4289 DVDD:5472 DVDD:5504 0.236776
rDVDD/4290 DVDD:5472 DVDD:5489 1.73333
rDVDD/4291 DVDD:5469 DVDD:5472 0.377206
rDVDD/4292 DVDD:5469 DVDD:5489 1.73333
rDVDD/4293 DVDD:5466 DVDD:5488 0.490893
rDVDD/4294 DVDD:5466 DVDD:5469 0.377206
rDVDD/4295 DVDD:5466 DVDD:5489 1.73333
rDVDD/4296 DVDD:5461 DVDD:5496 0.236794
rDVDD/4297 DVDD:5461 DVDD:5481 1.73333
rDVDD/4298 DVDD:5458 DVDD:5461 0.377206
rDVDD/4299 DVDD:5458 DVDD:5481 1.73333
rDVDD/4300 DVDD:5455 DVDD:5480 0.490911
rDVDD/4301 DVDD:5455 DVDD:5458 0.377206
rDVDD/4302 DVDD:5455 DVDD:5481 1.73333
rDVDD/4303 X49/X0/X2/X0/C0:pos DVDD:5481 3.65613
rDVDD/4304 X49/X0/X2/X0/C0:pos DVDD:5489 3.6566
rDVDD/4305 DVDD:5394 DVDD:12367 0.01368
rDVDD/4306 DVDD:5386 DVDD:12340 0.013662
rDVDD/4307 DVDD:5379 DVDD:5394 0.52
rDVDD/4308 DVDD:5378 DVDD:5379 0.433333
rDVDD/4309 DVDD:5371 DVDD:5386 0.52
rDVDD/4310 DVDD:5370 DVDD:5378 0.280062
rDVDD/4311 DVDD:5370 DVDD:5371 0.433333
rDVDD/4312 DVDD:5362 DVDD:5394 0.236776
rDVDD/4313 DVDD:5362 DVDD:5379 1.73333
rDVDD/4314 DVDD:5359 DVDD:5362 0.377206
rDVDD/4315 DVDD:5359 DVDD:5379 1.73333
rDVDD/4316 DVDD:5356 DVDD:5378 0.490893
rDVDD/4317 DVDD:5356 DVDD:5359 0.377206
rDVDD/4318 DVDD:5356 DVDD:5379 1.73333
rDVDD/4319 DVDD:5351 DVDD:5386 0.236794
rDVDD/4320 DVDD:5351 DVDD:5371 1.73333
rDVDD/4321 DVDD:5348 DVDD:5351 0.377206
rDVDD/4322 DVDD:5348 DVDD:5371 1.73333
rDVDD/4323 DVDD:5345 DVDD:5370 0.490911
rDVDD/4324 DVDD:5345 DVDD:5348 0.377206
rDVDD/4325 DVDD:5345 DVDD:5371 1.73333
rDVDD/4326 X49/X0/X1/X1/C0:pos DVDD:5371 3.65613
rDVDD/4327 X49/X0/X1/X1/C0:pos DVDD:5379 3.6566
rDVDD/4328 DVDD:5332 DVDD:11946 0.01368
rDVDD/4329 DVDD:5324 DVDD:11919 0.013662
rDVDD/4330 DVDD:5317 DVDD:5332 0.52
rDVDD/4331 DVDD:5316 DVDD:11188 0.0117
rDVDD/4332 DVDD:5316 DVDD:5317 0.433333
rDVDD/4333 DVDD:5309 DVDD:5324 0.52
rDVDD/4334 DVDD:5308 DVDD:11159 0.011682
rDVDD/4335 DVDD:5308 DVDD:5309 0.433333
rDVDD/4336 DVDD:5300 DVDD:5332 0.236776
rDVDD/4337 DVDD:5300 DVDD:5317 1.73333
rDVDD/4338 DVDD:5297 DVDD:5300 0.377206
rDVDD/4339 DVDD:5297 DVDD:5317 1.73333
rDVDD/4340 DVDD:5294 DVDD:5316 0.490893
rDVDD/4341 DVDD:5294 DVDD:5297 0.377206
rDVDD/4342 DVDD:5294 DVDD:5317 1.73333
rDVDD/4343 DVDD:5289 DVDD:5324 0.236794
rDVDD/4344 DVDD:5289 DVDD:5309 1.73333
rDVDD/4345 DVDD:5286 DVDD:5289 0.377206
rDVDD/4346 DVDD:5286 DVDD:5309 1.73333
rDVDD/4347 DVDD:5283 DVDD:5308 0.490911
rDVDD/4348 DVDD:5283 DVDD:5286 0.377206
rDVDD/4349 DVDD:5283 DVDD:5309 1.73333
rDVDD/4350 X49/X0/X1/X0/C0:pos DVDD:5309 3.65613
rDVDD/4351 X49/X0/X1/X0/C0:pos DVDD:5317 3.6566
rDVDD/4352 DVDD:5116 DVDD:13592 0.0117
rDVDD/4353 DVDD:5108 DVDD:13565 0.011682
rDVDD/4354 DVDD:5101 DVDD:5116 0.52
rDVDD/4355 DVDD:5100 DVDD:13277 0.01368
rDVDD/4356 DVDD:5100 DVDD:5101 0.433333
rDVDD/4357 DVDD:5093 DVDD:5108 0.52
rDVDD/4358 DVDD:5092 DVDD:13250 0.013662
rDVDD/4359 DVDD:5092 DVDD:5093 0.433333
rDVDD/4360 DVDD:5084 DVDD:5116 0.236776
rDVDD/4361 DVDD:5084 DVDD:5101 1.73333
rDVDD/4362 DVDD:5081 DVDD:5084 0.377206
rDVDD/4363 DVDD:5081 DVDD:5101 1.73333
rDVDD/4364 DVDD:5078 DVDD:5100 0.490893
rDVDD/4365 DVDD:5078 DVDD:5081 0.377206
rDVDD/4366 DVDD:5078 DVDD:5101 1.73333
rDVDD/4367 DVDD:5073 DVDD:5108 0.236794
rDVDD/4368 DVDD:5073 DVDD:5093 1.73333
rDVDD/4369 DVDD:5070 DVDD:5073 0.377206
rDVDD/4370 DVDD:5070 DVDD:5093 1.73333
rDVDD/4371 DVDD:5067 DVDD:5092 0.490911
rDVDD/4372 DVDD:5067 DVDD:5070 0.377206
rDVDD/4373 DVDD:5067 DVDD:5093 1.73333
rDVDD/4374 X48/X2/X1/C0:pos DVDD:5093 3.65613
rDVDD/4375 X48/X2/X1/C0:pos DVDD:5101 3.6566
rDVDD/4376 DVDD:5046 DVDD:5054 0.280062
rDVDD/4377 DVDD:5039 DVDD:5054 0.52
rDVDD/4378 DVDD:5038 DVDD:12962 0.01368
rDVDD/4379 DVDD:5038 DVDD:5039 0.433333
rDVDD/4380 DVDD:5031 DVDD:5046 0.52
rDVDD/4381 DVDD:5030 DVDD:12935 0.013662
rDVDD/4382 DVDD:5030 DVDD:5031 0.433333
rDVDD/4383 DVDD:5022 DVDD:5054 0.236776
rDVDD/4384 DVDD:5022 DVDD:5039 1.73333
rDVDD/4385 DVDD:5019 DVDD:5022 0.377206
rDVDD/4386 DVDD:5019 DVDD:5039 1.73333
rDVDD/4387 DVDD:5016 DVDD:5038 0.490893
rDVDD/4388 DVDD:5016 DVDD:5019 0.377206
rDVDD/4389 DVDD:5016 DVDD:5039 1.73333
rDVDD/4390 DVDD:5011 DVDD:5046 0.236794
rDVDD/4391 DVDD:5011 DVDD:5031 1.73333
rDVDD/4392 DVDD:5008 DVDD:5011 0.377206
rDVDD/4393 DVDD:5008 DVDD:5031 1.73333
rDVDD/4394 DVDD:5005 DVDD:5030 0.490911
rDVDD/4395 DVDD:5005 DVDD:5008 0.377206
rDVDD/4396 DVDD:5005 DVDD:5031 1.73333
rDVDD/4397 X48/X2/X0/C0:pos DVDD:5031 3.65613
rDVDD/4398 X48/X2/X0/C0:pos DVDD:5039 3.6566
rDVDD/4399 DVDD:4944 DVDD:12647 0.01368
rDVDD/4400 DVDD:4936 DVDD:12620 0.013662
rDVDD/4401 DVDD:4929 DVDD:4944 0.52
rDVDD/4402 DVDD:4928 DVDD:4929 0.433333
rDVDD/4403 DVDD:4921 DVDD:4936 0.52
rDVDD/4404 DVDD:4920 DVDD:4928 0.280062
rDVDD/4405 DVDD:4920 DVDD:4921 0.433333
rDVDD/4406 DVDD:4912 DVDD:4944 0.236776
rDVDD/4407 DVDD:4912 DVDD:4929 1.73333
rDVDD/4408 DVDD:4909 DVDD:4912 0.377206
rDVDD/4409 DVDD:4909 DVDD:4929 1.73333
rDVDD/4410 DVDD:4906 DVDD:4928 0.490893
rDVDD/4411 DVDD:4906 DVDD:4909 0.377206
rDVDD/4412 DVDD:4906 DVDD:4929 1.73333
rDVDD/4413 DVDD:4901 DVDD:4936 0.236794
rDVDD/4414 DVDD:4901 DVDD:4921 1.73333
rDVDD/4415 DVDD:4898 DVDD:4901 0.377206
rDVDD/4416 DVDD:4898 DVDD:4921 1.73333
rDVDD/4417 DVDD:4895 DVDD:4920 0.490911
rDVDD/4418 DVDD:4895 DVDD:4898 0.377206
rDVDD/4419 DVDD:4895 DVDD:4921 1.73333
rDVDD/4420 X48/X1/X1/C0:pos DVDD:4921 3.65613
rDVDD/4421 X48/X1/X1/C0:pos DVDD:4929 3.6566
rDVDD/4422 DVDD:4882 DVDD:12226 0.01368
rDVDD/4423 DVDD:4874 DVDD:12199 0.013662
rDVDD/4424 DVDD:4867 DVDD:4882 0.52
rDVDD/4425 DVDD:4866 DVDD:10734 0.0117
rDVDD/4426 DVDD:4866 DVDD:4867 0.433333
rDVDD/4427 DVDD:4859 DVDD:4874 0.52
rDVDD/4428 DVDD:4858 DVDD:10772 0.000522
rDVDD/4429 DVDD:4858 DVDD:4859 0.433333
rDVDD/4430 DVDD:4850 DVDD:4882 0.236776
rDVDD/4431 DVDD:4850 DVDD:4867 1.73333
rDVDD/4432 DVDD:4847 DVDD:4850 0.377206
rDVDD/4433 DVDD:4847 DVDD:4867 1.73333
rDVDD/4434 DVDD:4844 DVDD:4866 0.490893
rDVDD/4435 DVDD:4844 DVDD:4847 0.377206
rDVDD/4436 DVDD:4844 DVDD:4867 1.73333
rDVDD/4437 DVDD:4839 DVDD:4874 0.236794
rDVDD/4438 DVDD:4839 DVDD:4859 1.73333
rDVDD/4439 DVDD:4836 DVDD:4839 0.377206
rDVDD/4440 DVDD:4836 DVDD:4859 1.73333
rDVDD/4441 DVDD:4833 DVDD:4858 0.490911
rDVDD/4442 DVDD:4833 DVDD:4836 0.377206
rDVDD/4443 DVDD:4833 DVDD:4859 1.73333
rDVDD/4444 X48/X1/X0/C0:pos DVDD:4859 3.65613
rDVDD/4445 X48/X1/X0/C0:pos DVDD:4867 3.6566
rDVDD/4446 DVDD:4225 DVDD:15249 0.464528
rDVDD/4447 DVDD:4225 DVDD:4226 0.28125
rDVDD/4448 DVDD:4223 DVDD:15261 0.0552756
rDVDD/4449 DVDD:4223 DVDD:15265 0.0325984
rDVDD/4450 DVDD:4223 DVDD:4224 0.28125
rDVDD/4451 DVDD:4221 DVDD:4222 1.125
rDVDD/4452 DVDD:4219 DVDD:4221 0.0382677
rDVDD/4453 DVDD:4219 DVDD:4220 1.125
rDVDD/4454 DVDD:4217 DVDD:4219 0.0382677
rDVDD/4455 DVDD:4217 DVDD:4218 1.125
rDVDD/4456 DVDD:4215 DVDD:4217 0.0382677
rDVDD/4457 DVDD:4215 DVDD:4216 1.125
rDVDD/4458 DVDD:4213 DVDD:4215 0.0382677
rDVDD/4459 DVDD:4211 DVDD:4212 1.125
rDVDD/4460 DVDD:4209 DVDD:4211 0.0382677
rDVDD/4461 DVDD:4209 DVDD:4210 1.125
rDVDD/4462 DVDD:4207 DVDD:4209 0.0382677
rDVDD/4463 DVDD:4207 DVDD:4208 1.125
rDVDD/4464 DVDD:4205 DVDD:4207 0.0382677
rDVDD/4465 DVDD:4205 DVDD:4206 1.125
rDVDD/4466 DVDD:4203 DVDD:4205 0.0382677
rDVDD/4467 DVDD:4201 DVDD:4202 1.125
rDVDD/4468 DVDD:4199 DVDD:4201 0.0382677
rDVDD/4469 DVDD:4199 DVDD:4200 1.125
rDVDD/4470 DVDD:4197 DVDD:4199 0.0382677
rDVDD/4471 DVDD:4197 DVDD:4198 1.125
rDVDD/4472 DVDD:4195 DVDD:4197 0.0382677
rDVDD/4473 DVDD:4195 DVDD:4196 1.125
rDVDD/4474 DVDD:4193 DVDD:4195 0.0382677
rDVDD/4475 DVDD:4193 DVDD:4194 2.25
rDVDD/4476 DVDD:4191 DVDD:4192 1.125
rDVDD/4477 DVDD:4189 DVDD:4191 0.0382677
rDVDD/4478 DVDD:4189 DVDD:4190 1.125
rDVDD/4479 DVDD:4187 DVDD:4189 0.0382677
rDVDD/4480 DVDD:4187 DVDD:4188 1.125
rDVDD/4481 DVDD:4185 DVDD:4187 0.0382677
rDVDD/4482 DVDD:4185 DVDD:4186 1.125
rDVDD/4483 DVDD:4183 DVDD:4185 0.0382677
rDVDD/4484 DVDD:4182 DVDD:4222 0.058386
rDVDD/4485 DVDD:4182 DVDD:4221 1.16327
rDVDD/4486 DVDD:4179 DVDD:4213 0.0191339
rDVDD/4487 DVDD:4178 DVDD:4179 1.125
rDVDD/4488 DVDD:4178 DVDD:4212 0.0908548
rDVDD/4489 DVDD:4177 DVDD:4179 0.0382677
rDVDD/4490 DVDD:4177 DVDD:4211 0.0382677
rDVDD/4491 DVDD:4177 DVDD:4178 1.125
rDVDD/4492 DVDD:4175 DVDD:4203 0.0191339
rDVDD/4493 DVDD:4174 DVDD:4175 1.125
rDVDD/4494 DVDD:4174 DVDD:4202 0.0908548
rDVDD/4495 DVDD:4173 DVDD:4175 0.0382677
rDVDD/4496 DVDD:4173 DVDD:4201 0.0382677
rDVDD/4497 DVDD:4173 DVDD:4174 1.125
rDVDD/4498 DVDD:4171 DVDD:4193 0.0191339
rDVDD/4499 DVDD:4170 DVDD:4194 0.0908548
rDVDD/4500 DVDD:4170 DVDD:4171 1.125
rDVDD/4501 DVDD:4170 DVDD:4192 0.0908548
rDVDD/4502 DVDD:4169 DVDD:4171 0.0382677
rDVDD/4503 DVDD:4169 DVDD:4191 0.0382677
rDVDD/4504 DVDD:4169 DVDD:4170 1.125
rDVDD/4505 DVDD:4167 DVDD:4183 0.0191339
rDVDD/4506 DVDD:4167 DVDD:4225 0.256713
rDVDD/4507 DVDD:4167 DVDD:4168 1.125
rDVDD/4508 DVDD:4165 DVDD:4166 1.5
rDVDD/4509 DVDD:4163 DVDD:4164 1.5
rDVDD/4510 DVDD:4161 DVDD:4165 0.0191339
rDVDD/4511 DVDD:4159 DVDD:4161 0.225531
rDVDD/4512 DVDD:4159 DVDD:4160 0.5625
rDVDD/4513 DVDD:4157 DVDD:4159 0.24874
rDVDD/4514 DVDD:4157 DVDD:4158 0.5625
rDVDD/4515 DVDD:4155 DVDD:4157 0.24874
rDVDD/4516 DVDD:4155 DVDD:4163 0.225531
rDVDD/4517 DVDD:4155 DVDD:4156 0.5625
rDVDD/4518 DVDD:4153 DVDD:4163 0.0191339
rDVDD/4519 DVDD:4151 DVDD:4153 0.232087
rDVDD/4520 DVDD:4151 DVDD:14949 0.464528
rDVDD/4521 DVDD:4151 DVDD:4152 0.28125
rDVDD/4522 DVDD:4149 DVDD:14961 0.0333071
rDVDD/4523 DVDD:4149 DVDD:14965 0.0545669
rDVDD/4524 DVDD:4149 DVDD:4150 0.28125
rDVDD/4525 DVDD:4148 DVDD:4165 1.5
rDVDD/4526 DVDD:4146 DVDD:4159 0.642857
rDVDD/4527 DVDD:4144 DVDD:4157 0.642857
rDVDD/4528 DVDD:4142 DVDD:4155 0.642857
rDVDD/4529 DVDD:4140 DVDD:4163 1.5
rDVDD/4530 DVDD:4138 DVDD:4161 4.5
rDVDD/4531 DVDD:4138 DVDD:4148 0.0437838
rDVDD/4532 DVDD:4136 DVDD:4153 4.5
rDVDD/4533 DVDD:4136 DVDD:4140 0.0437838
rDVDD/4534 DVDD:4133 DVDD:4134 1.5
rDVDD/4535 DVDD:4131 DVDD:4132 1.5
rDVDD/4536 DVDD:4129 DVDD:4133 0.0191339
rDVDD/4537 DVDD:4127 DVDD:4129 0.225531
rDVDD/4538 DVDD:4127 DVDD:4128 0.5625
rDVDD/4539 DVDD:4125 DVDD:4127 0.24874
rDVDD/4540 DVDD:4125 DVDD:4126 0.5625
rDVDD/4541 DVDD:4123 DVDD:4125 0.24874
rDVDD/4542 DVDD:4123 DVDD:4131 0.225531
rDVDD/4543 DVDD:4123 DVDD:4124 0.5625
rDVDD/4544 DVDD:4121 DVDD:4131 0.0191339
rDVDD/4545 DVDD:4119 DVDD:4121 0.232087
rDVDD/4546 DVDD:4119 DVDD:14664 0.464528
rDVDD/4547 DVDD:4119 DVDD:4120 0.28125
rDVDD/4548 DVDD:4117 DVDD:14676 0.0552756
rDVDD/4549 DVDD:4117 DVDD:14680 0.0325984
rDVDD/4550 DVDD:4117 DVDD:4118 0.28125
rDVDD/4551 DVDD:4116 DVDD:4133 1.5
rDVDD/4552 DVDD:4114 DVDD:4127 0.642857
rDVDD/4553 DVDD:4112 DVDD:4125 0.642857
rDVDD/4554 DVDD:4110 DVDD:4123 0.642857
rDVDD/4555 DVDD:4108 DVDD:4131 1.5
rDVDD/4556 DVDD:4106 DVDD:4129 4.5
rDVDD/4557 DVDD:4104 DVDD:4121 4.5
rDVDD/4558 DVDD:4101 DVDD:4102 1.5
rDVDD/4559 DVDD:4099 DVDD:4100 1.5
rDVDD/4560 DVDD:4098 DVDD:4102 0.0437838
rDVDD/4561 DVDD:4097 DVDD:4101 0.0191339
rDVDD/4562 DVDD:4097 DVDD:4098 1.5
rDVDD/4563 DVDD:4095 DVDD:4097 0.225531
rDVDD/4564 DVDD:4093 DVDD:4095 0.24874
rDVDD/4565 DVDD:4091 DVDD:4093 0.24874
rDVDD/4566 DVDD:4091 DVDD:4099 0.225531
rDVDD/4567 DVDD:4090 DVDD:4100 0.0437838
rDVDD/4568 DVDD:4089 DVDD:4099 0.0191339
rDVDD/4569 DVDD:4089 DVDD:4090 1.5
rDVDD/4570 DVDD:4087 DVDD:4089 0.232087
rDVDD/4571 DVDD:4087 DVDD:14379 0.464528
rDVDD/4572 DVDD:4087 DVDD:4088 0.28125
rDVDD/4573 DVDD:4085 DVDD:14391 0.0552756
rDVDD/4574 DVDD:4085 DVDD:14395 0.0325984
rDVDD/4575 DVDD:4085 DVDD:4086 0.28125
rDVDD/4576 DVDD:4084 DVDD:4101 1.5
rDVDD/4577 DVDD:4082 DVDD:4095 0.642857
rDVDD/4578 DVDD:4080 DVDD:4093 0.642857
rDVDD/4579 DVDD:4078 DVDD:4091 0.642857
rDVDD/4580 DVDD:4076 DVDD:4099 1.5
rDVDD/4581 DVDD:4074 DVDD:4097 4.5
rDVDD/4582 DVDD:4074 DVDD:4084 0.0437838
rDVDD/4583 DVDD:4072 DVDD:4089 4.5
rDVDD/4584 DVDD:4072 DVDD:4076 0.0437838
rDVDD/4585 DVDD:4069 DVDD:4070 1.5
rDVDD/4586 DVDD:4067 DVDD:4068 1.5
rDVDD/4587 DVDD:4066 DVDD:4070 0.0437838
rDVDD/4588 DVDD:4065 DVDD:4069 0.0191339
rDVDD/4589 DVDD:4065 DVDD:4066 1.5
rDVDD/4590 DVDD:4063 DVDD:4065 0.225531
rDVDD/4591 DVDD:4063 DVDD:4064 0.5625
rDVDD/4592 DVDD:4061 DVDD:4063 0.24874
rDVDD/4593 DVDD:4061 DVDD:4062 0.5625
rDVDD/4594 DVDD:4059 DVDD:4061 0.24874
rDVDD/4595 DVDD:4059 DVDD:4067 0.225531
rDVDD/4596 DVDD:4059 DVDD:4060 0.5625
rDVDD/4597 DVDD:4058 DVDD:4068 0.0437838
rDVDD/4598 DVDD:4057 DVDD:4067 0.0191339
rDVDD/4599 DVDD:4057 DVDD:4058 1.5
rDVDD/4600 DVDD:4055 DVDD:4057 0.232087
rDVDD/4601 DVDD:4055 DVDD:14100 0.464528
rDVDD/4602 DVDD:4055 DVDD:4056 0.28125
rDVDD/4603 DVDD:4053 DVDD:14112 0.0333071
rDVDD/4604 DVDD:4053 DVDD:14116 0.0545669
rDVDD/4605 DVDD:4053 DVDD:4054 0.28125
rDVDD/4606 DVDD:4052 DVDD:4069 1.5
rDVDD/4607 DVDD:4050 DVDD:4063 0.642857
rDVDD/4608 DVDD:4048 DVDD:4061 0.642857
rDVDD/4609 DVDD:4046 DVDD:4059 0.642857
rDVDD/4610 DVDD:4044 DVDD:4067 1.5
rDVDD/4611 DVDD:4042 DVDD:4065 4.5
rDVDD/4612 DVDD:4042 DVDD:4052 0.0437838
rDVDD/4613 DVDD:4040 DVDD:4057 4.5
rDVDD/4614 DVDD:4040 DVDD:4044 0.0437838
rDVDD/4615 DVDD:4037 DVDD:13915 0.464528
rDVDD/4616 DVDD:4037 DVDD:4038 0.28125
rDVDD/4617 DVDD:4035 DVDD:13927 0.0552756
rDVDD/4618 DVDD:4035 DVDD:13931 0.0325984
rDVDD/4619 DVDD:4035 DVDD:4036 0.28125
rDVDD/4620 DVDD:4033 DVDD:4034 1.125
rDVDD/4621 DVDD:4031 DVDD:4033 0.0382677
rDVDD/4622 DVDD:4031 DVDD:4032 1.125
rDVDD/4623 DVDD:4029 DVDD:4031 0.0382677
rDVDD/4624 DVDD:4029 DVDD:4030 1.125
rDVDD/4625 DVDD:4027 DVDD:4029 0.0382677
rDVDD/4626 DVDD:4027 DVDD:4028 1.125
rDVDD/4627 DVDD:4025 DVDD:4027 0.0382677
rDVDD/4628 DVDD:4025 DVDD:4026 2.25
rDVDD/4629 DVDD:4023 DVDD:4024 1.125
rDVDD/4630 DVDD:4021 DVDD:4023 0.0382677
rDVDD/4631 DVDD:4021 DVDD:4022 1.125
rDVDD/4632 DVDD:4019 DVDD:4021 0.0382677
rDVDD/4633 DVDD:4019 DVDD:4020 1.125
rDVDD/4634 DVDD:4017 DVDD:4019 0.0382677
rDVDD/4635 DVDD:4017 DVDD:4018 1.125
rDVDD/4636 DVDD:4015 DVDD:4017 0.0382677
rDVDD/4637 DVDD:4015 DVDD:4016 2.25
rDVDD/4638 DVDD:4013 DVDD:4014 1.125
rDVDD/4639 DVDD:4011 DVDD:4013 0.0382677
rDVDD/4640 DVDD:4011 DVDD:4012 1.125
rDVDD/4641 DVDD:4009 DVDD:4011 0.0382677
rDVDD/4642 DVDD:4009 DVDD:4010 1.125
rDVDD/4643 DVDD:4007 DVDD:4009 0.0382677
rDVDD/4644 DVDD:4007 DVDD:4008 1.125
rDVDD/4645 DVDD:4005 DVDD:4007 0.0382677
rDVDD/4646 DVDD:4005 DVDD:4006 2.25
rDVDD/4647 DVDD:4003 DVDD:4004 1.125
rDVDD/4648 DVDD:4001 DVDD:4003 0.0382677
rDVDD/4649 DVDD:4001 DVDD:4002 1.125
rDVDD/4650 DVDD:3999 DVDD:4001 0.0382677
rDVDD/4651 DVDD:3999 DVDD:4000 1.125
rDVDD/4652 DVDD:3997 DVDD:3999 0.0382677
rDVDD/4653 DVDD:3997 DVDD:3998 1.125
rDVDD/4654 DVDD:3995 DVDD:3997 0.0382677
rDVDD/4655 DVDD:3994 DVDD:4034 0.058386
rDVDD/4656 DVDD:3994 DVDD:4033 1.16327
rDVDD/4657 DVDD:3991 DVDD:4025 0.0191339
rDVDD/4658 DVDD:3990 DVDD:4026 0.0908548
rDVDD/4659 DVDD:3990 DVDD:3991 1.125
rDVDD/4660 DVDD:3990 DVDD:4024 0.0908548
rDVDD/4661 DVDD:3989 DVDD:3991 0.0382677
rDVDD/4662 DVDD:3989 DVDD:4023 0.0382677
rDVDD/4663 DVDD:3989 DVDD:3990 1.125
rDVDD/4664 DVDD:3987 DVDD:4015 0.0191339
rDVDD/4665 DVDD:3986 DVDD:4016 0.0908548
rDVDD/4666 DVDD:3986 DVDD:3987 1.125
rDVDD/4667 DVDD:3986 DVDD:4014 0.0908548
rDVDD/4668 DVDD:3985 DVDD:3987 0.0382677
rDVDD/4669 DVDD:3985 DVDD:4013 0.0382677
rDVDD/4670 DVDD:3985 DVDD:3986 1.125
rDVDD/4671 DVDD:3983 DVDD:4005 0.0191339
rDVDD/4672 DVDD:3982 DVDD:4006 0.0908548
rDVDD/4673 DVDD:3982 DVDD:3983 1.125
rDVDD/4674 DVDD:3982 DVDD:4004 0.0908548
rDVDD/4675 DVDD:3981 DVDD:3983 0.0382677
rDVDD/4676 DVDD:3981 DVDD:4003 0.0382677
rDVDD/4677 DVDD:3981 DVDD:3982 1.125
rDVDD/4678 DVDD:3979 DVDD:3995 0.0191339
rDVDD/4679 DVDD:3979 DVDD:4037 0.256713
rDVDD/4680 DVDD:3979 DVDD:3980 1.125
rDVDD/4681 DVDD:2246 DVDD:4036 0.0238077
rDVDD/4682 DVDD:2246 X46/D0:neg 0.709092
rDVDD/4683 DVDD:2244 DVDD:4036 0.0146538
rDVDD/4684 DVDD:2244 X46/D0:neg 0.709092
rDVDD/4685 DVDD:2242 DVDD:2244 0.0384615
rDVDD/4686 DVDD:2242 X46/D0:neg 0.354546
rDVDD/4687 DVDD:2238 DVDD:2242 0.0384615
rDVDD/4688 DVDD:2238 X46/D0:neg 0.709092
rDVDD/4689 DVDD:2236 DVDD:2238 0.0384615
rDVDD/4690 DVDD:2236 X46/D0:neg 0.354546
rDVDD/4691 DVDD:2232 DVDD:2236 0.0384615
rDVDD/4692 DVDD:2232 X46/D0:neg 0.709092
rDVDD/4693 DVDD:2230 DVDD:2232 0.0576923
rDVDD/4694 DVDD:2230 X46/D0:neg 0.354546
rDVDD/4695 DVDD:2226 DVDD:2230 0.0384615
rDVDD/4696 DVDD:2226 X46/D0:neg 0.709092
rDVDD/4697 DVDD:2224 DVDD:2226 0.0384615
rDVDD/4698 DVDD:2224 DVDD:4054 0.0245769
rDVDD/4699 DVDD:2224 X46/D0:neg 0.354546
rDVDD/4700 DVDD:2220 DVDD:4054 0.0138846
rDVDD/4701 DVDD:2220 X46/D0:neg 0.709092
rDVDD/4702 DVDD:2218 DVDD:2220 0.0384615
rDVDD/4703 DVDD:2218 X46/D0:neg 0.709092
rDVDD/4704 DVDD:2216 DVDD:2218 0.0192308
rDVDD/4705 DVDD:2216 X46/D0:neg 0.709092
rDVDD/4706 DVDD:2214 DVDD:2216 0.0384615
rDVDD/4707 DVDD:2214 X46/D0:neg 0.709092
rDVDD/4708 DVDD:2212 DVDD:2214 0.0384615
rDVDD/4709 DVDD:2212 X46/D0:neg 0.354546
rDVDD/4710 DVDD:2208 DVDD:2212 0.0384615
rDVDD/4711 DVDD:2208 X46/D0:neg 0.709092
rDVDD/4712 DVDD:2206 DVDD:2208 0.0384615
rDVDD/4713 DVDD:2206 X46/D0:neg 0.354546
rDVDD/4714 DVDD:2202 DVDD:2206 0.0384615
rDVDD/4715 DVDD:2202 X46/D0:neg 0.709092
rDVDD/4716 DVDD:2200 DVDD:2202 0.0576923
rDVDD/4717 DVDD:2200 X46/D0:neg 0.354546
rDVDD/4718 DVDD:2196 DVDD:2200 0.0384615
rDVDD/4719 DVDD:2196 X46/D0:neg 0.709092
rDVDD/4720 DVDD:2194 DVDD:2196 0.0384615
rDVDD/4721 DVDD:2194 DVDD:4086 0.0384231
rDVDD/4722 DVDD:2194 X46/D0:neg 0.354546
rDVDD/4723 DVDD:2190 DVDD:4086 3.84615e-05
rDVDD/4724 DVDD:2190 X46/D0:neg 0.709092
rDVDD/4725 DVDD:2188 DVDD:2190 0.0384615
rDVDD/4726 DVDD:2188 X46/D0:neg 0.709092
rDVDD/4727 DVDD:2186 DVDD:2188 0.0192308
rDVDD/4728 DVDD:2186 X46/D0:neg 0.709092
rDVDD/4729 DVDD:2184 DVDD:2186 0.0384615
rDVDD/4730 DVDD:2184 X46/D0:neg 0.709092
rDVDD/4731 DVDD:2182 DVDD:2184 0.0384615
rDVDD/4732 DVDD:2182 X46/D0:neg 0.354546
rDVDD/4733 DVDD:2178 DVDD:2182 0.0384615
rDVDD/4734 DVDD:2178 X46/D0:neg 0.709092
rDVDD/4735 DVDD:2176 DVDD:2178 0.0384615
rDVDD/4736 DVDD:2176 X46/D0:neg 0.354546
rDVDD/4737 DVDD:2172 DVDD:2176 0.0384615
rDVDD/4738 DVDD:2172 X46/D0:neg 0.709092
rDVDD/4739 DVDD:2170 DVDD:2172 0.0576538
rDVDD/4740 DVDD:2170 X46/D0:neg 0.354546
rDVDD/4741 DVDD:2166 DVDD:2170 0.0384615
rDVDD/4742 DVDD:2166 X46/D0:neg 0.709092
rDVDD/4743 DVDD:2164 DVDD:2166 0.0384615
rDVDD/4744 DVDD:2164 X46/D0:neg 0.354546
rDVDD/4745 DVDD:2160 DVDD:2164 0.0384615
rDVDD/4746 DVDD:2160 X46/D0:neg 0.709092
rDVDD/4747 DVDD:2158 DVDD:2160 0.0384615
rDVDD/4748 DVDD:2158 X46/D0:neg 0.709092
rDVDD/4749 DVDD:2156 DVDD:2158 0.0192308
rDVDD/4750 DVDD:2156 DVDD:4118 0.0338462
rDVDD/4751 DVDD:2156 X46/D0:neg 0.709092
rDVDD/4752 DVDD:2154 DVDD:4118 0.00461538
rDVDD/4753 DVDD:2154 X46/D0:neg 0.709092
rDVDD/4754 DVDD:2152 DVDD:2154 0.0384615
rDVDD/4755 DVDD:2152 X46/D0:neg 0.354546
rDVDD/4756 DVDD:2148 DVDD:2152 0.0384615
rDVDD/4757 DVDD:2148 X46/D0:neg 0.709092
rDVDD/4758 DVDD:2146 DVDD:2148 0.0384615
rDVDD/4759 DVDD:2146 X46/D0:neg 0.354546
rDVDD/4760 DVDD:2142 DVDD:2146 0.0384615
rDVDD/4761 DVDD:2142 X46/D0:neg 0.709092
rDVDD/4762 DVDD:2140 DVDD:2142 0.0576923
rDVDD/4763 DVDD:2140 X46/D0:neg 0.354546
rDVDD/4764 DVDD:2136 DVDD:2140 0.0384615
rDVDD/4765 DVDD:2136 X46/D0:neg 0.709092
rDVDD/4766 DVDD:2134 DVDD:2136 0.0384615
rDVDD/4767 DVDD:2134 X46/D0:neg 0.354546
rDVDD/4768 DVDD:2130 DVDD:2134 0.0384615
rDVDD/4769 DVDD:2130 X46/D0:neg 0.709092
rDVDD/4770 DVDD:2128 DVDD:2130 0.0384615
rDVDD/4771 DVDD:2128 X46/D0:neg 0.709092
rDVDD/4772 DVDD:2126 DVDD:2128 0.0192308
rDVDD/4773 DVDD:2126 X46/D0:neg 0.709092
rDVDD/4774 DVDD:2124 DVDD:2126 0.0384615
rDVDD/4775 DVDD:2124 DVDD:4150 0.00923077
rDVDD/4776 DVDD:2124 X46/D0:neg 0.709092
rDVDD/4777 DVDD:2122 DVDD:4150 0.0292308
rDVDD/4778 DVDD:2122 X46/D0:neg 0.354546
rDVDD/4779 DVDD:2118 DVDD:2122 0.0384615
rDVDD/4780 DVDD:2118 X46/D0:neg 0.709092
rDVDD/4781 DVDD:2116 DVDD:2118 0.0384615
rDVDD/4782 DVDD:2116 X46/D0:neg 0.354546
rDVDD/4783 DVDD:2112 DVDD:2116 0.0384615
rDVDD/4784 DVDD:2112 X46/D0:neg 0.709092
rDVDD/4785 DVDD:2110 DVDD:2112 0.0576923
rDVDD/4786 DVDD:2110 X46/D0:neg 0.354546
rDVDD/4787 DVDD:2106 DVDD:2110 0.0384615
rDVDD/4788 DVDD:2106 X46/D0:neg 0.709092
rDVDD/4789 DVDD:2104 DVDD:2106 0.0384615
rDVDD/4790 DVDD:2104 X46/D0:neg 0.354546
rDVDD/4791 DVDD:2100 DVDD:2104 0.0384615
rDVDD/4792 DVDD:2100 DVDD:4224 0.01
rDVDD/4793 DVDD:2100 X46/D0:neg 0.709092
rDVDD/4794 DVDD:2098 DVDD:4224 0.0284615
rDVDD/4795 DVDD:2098 X46/D0:neg 0.709092
rDVDD/4796 DVDD:2096 DVDD:2098 0.0192308
rDVDD/4797 DVDD:2096 X46/D0:neg 1.04
rDVDD/4798 DVDD:2093 DVDD:4038 0.0238077
rDVDD/4799 DVDD:2093 X46/D0:neg 0.709092
rDVDD/4800 DVDD:2091 DVDD:4038 0.0146538
rDVDD/4801 DVDD:2091 X46/D0:neg 0.709092
rDVDD/4802 DVDD:2089 DVDD:2091 0.0384615
rDVDD/4803 DVDD:2089 X46/D0:neg 0.354546
rDVDD/4804 DVDD:2085 DVDD:2089 0.0384615
rDVDD/4805 DVDD:2085 X46/D0:neg 0.709092
rDVDD/4806 DVDD:2083 DVDD:2085 0.0384615
rDVDD/4807 DVDD:2083 X46/D0:neg 0.354546
rDVDD/4808 DVDD:2079 DVDD:2083 0.0384615
rDVDD/4809 DVDD:2079 X46/D0:neg 0.709092
rDVDD/4810 DVDD:2077 DVDD:2079 0.0576923
rDVDD/4811 DVDD:2077 X46/D0:neg 0.354546
rDVDD/4812 DVDD:2073 DVDD:2077 0.0384615
rDVDD/4813 DVDD:2073 X46/D0:neg 0.709092
rDVDD/4814 DVDD:2071 DVDD:2073 0.0384615
rDVDD/4815 DVDD:2071 DVDD:4056 0.0245769
rDVDD/4816 DVDD:2071 X46/D0:neg 0.354546
rDVDD/4817 DVDD:2067 DVDD:4056 0.0138846
rDVDD/4818 DVDD:2067 X46/D0:neg 0.709092
rDVDD/4819 DVDD:2065 DVDD:2067 0.0384615
rDVDD/4820 DVDD:2065 X46/D0:neg 0.709092
rDVDD/4821 DVDD:2063 DVDD:2065 0.0192308
rDVDD/4822 DVDD:2063 X46/D0:neg 0.709092
rDVDD/4823 DVDD:2061 DVDD:2063 0.0384615
rDVDD/4824 DVDD:2061 X46/D0:neg 0.709092
rDVDD/4825 DVDD:2059 DVDD:2061 0.0384615
rDVDD/4826 DVDD:2059 X46/D0:neg 0.354546
rDVDD/4827 DVDD:2055 DVDD:2059 0.0384615
rDVDD/4828 DVDD:2055 X46/D0:neg 0.709092
rDVDD/4829 DVDD:2053 DVDD:2055 0.0384615
rDVDD/4830 DVDD:2053 X46/D0:neg 0.354546
rDVDD/4831 DVDD:2049 DVDD:2053 0.0384615
rDVDD/4832 DVDD:2049 X46/D0:neg 0.709092
rDVDD/4833 DVDD:2047 DVDD:2049 0.0576923
rDVDD/4834 DVDD:2047 X46/D0:neg 0.354546
rDVDD/4835 DVDD:2043 DVDD:2047 0.0384615
rDVDD/4836 DVDD:2043 X46/D0:neg 0.709092
rDVDD/4837 DVDD:2041 DVDD:2043 0.0384615
rDVDD/4838 DVDD:2041 DVDD:4088 0.0384231
rDVDD/4839 DVDD:2041 X46/D0:neg 0.354546
rDVDD/4840 DVDD:2037 DVDD:4088 3.84615e-05
rDVDD/4841 DVDD:2037 X46/D0:neg 0.709092
rDVDD/4842 DVDD:2035 DVDD:2037 0.0384615
rDVDD/4843 DVDD:2035 X46/D0:neg 0.709092
rDVDD/4844 DVDD:2033 DVDD:2035 0.0192308
rDVDD/4845 DVDD:2033 X46/D0:neg 0.709092
rDVDD/4846 DVDD:2031 DVDD:2033 0.0384615
rDVDD/4847 DVDD:2031 X46/D0:neg 0.709092
rDVDD/4848 DVDD:2029 DVDD:2031 0.0384615
rDVDD/4849 DVDD:2029 X46/D0:neg 0.354546
rDVDD/4850 DVDD:2025 DVDD:2029 0.0384615
rDVDD/4851 DVDD:2025 X46/D0:neg 0.709092
rDVDD/4852 DVDD:2023 DVDD:2025 0.0384615
rDVDD/4853 DVDD:2023 X46/D0:neg 0.354546
rDVDD/4854 DVDD:2019 DVDD:2023 0.0384615
rDVDD/4855 DVDD:2019 X46/D0:neg 0.709092
rDVDD/4856 DVDD:2017 DVDD:2019 0.0576538
rDVDD/4857 DVDD:2017 X46/D0:neg 0.354546
rDVDD/4858 DVDD:2013 DVDD:2017 0.0384615
rDVDD/4859 DVDD:2013 X46/D0:neg 0.709092
rDVDD/4860 DVDD:2011 DVDD:2013 0.0384615
rDVDD/4861 DVDD:2011 X46/D0:neg 0.354546
rDVDD/4862 DVDD:2007 DVDD:2011 0.0384615
rDVDD/4863 DVDD:2007 X46/D0:neg 0.709092
rDVDD/4864 DVDD:2005 DVDD:2007 0.0384615
rDVDD/4865 DVDD:2005 X46/D0:neg 0.709092
rDVDD/4866 DVDD:2003 DVDD:2005 0.0192308
rDVDD/4867 DVDD:2003 DVDD:4120 0.0338462
rDVDD/4868 DVDD:2003 X46/D0:neg 0.709092
rDVDD/4869 DVDD:2001 DVDD:4120 0.00461538
rDVDD/4870 DVDD:2001 X46/D0:neg 0.709092
rDVDD/4871 DVDD:1999 DVDD:2001 0.0384615
rDVDD/4872 DVDD:1999 X46/D0:neg 0.354546
rDVDD/4873 DVDD:1995 DVDD:1999 0.0384615
rDVDD/4874 DVDD:1995 X46/D0:neg 0.709092
rDVDD/4875 DVDD:1993 DVDD:1995 0.0384615
rDVDD/4876 DVDD:1993 X46/D0:neg 0.354546
rDVDD/4877 DVDD:1989 DVDD:1993 0.0384615
rDVDD/4878 DVDD:1989 X46/D0:neg 0.709092
rDVDD/4879 DVDD:1987 DVDD:1989 0.0576923
rDVDD/4880 DVDD:1987 X46/D0:neg 0.354546
rDVDD/4881 DVDD:1983 DVDD:1987 0.0384615
rDVDD/4882 DVDD:1983 X46/D0:neg 0.709092
rDVDD/4883 DVDD:1981 DVDD:1983 0.0384615
rDVDD/4884 DVDD:1981 X46/D0:neg 0.354546
rDVDD/4885 DVDD:1977 DVDD:1981 0.0384615
rDVDD/4886 DVDD:1977 X46/D0:neg 0.709092
rDVDD/4887 DVDD:1975 DVDD:1977 0.0384615
rDVDD/4888 DVDD:1975 X46/D0:neg 0.709092
rDVDD/4889 DVDD:1973 DVDD:1975 0.0192308
rDVDD/4890 DVDD:1973 X46/D0:neg 0.709092
rDVDD/4891 DVDD:1971 DVDD:1973 0.0384615
rDVDD/4892 DVDD:1971 DVDD:4152 0.00923077
rDVDD/4893 DVDD:1971 X46/D0:neg 0.709092
rDVDD/4894 DVDD:1969 DVDD:4152 0.0292308
rDVDD/4895 DVDD:1969 X46/D0:neg 0.354546
rDVDD/4896 DVDD:1965 DVDD:1969 0.0384615
rDVDD/4897 DVDD:1965 X46/D0:neg 0.709092
rDVDD/4898 DVDD:1963 DVDD:1965 0.0384615
rDVDD/4899 DVDD:1963 X46/D0:neg 0.354546
rDVDD/4900 DVDD:1959 DVDD:1963 0.0384615
rDVDD/4901 DVDD:1959 X46/D0:neg 0.709092
rDVDD/4902 DVDD:1957 DVDD:1959 0.0576923
rDVDD/4903 DVDD:1957 X46/D0:neg 0.354546
rDVDD/4904 DVDD:1953 DVDD:1957 0.0384615
rDVDD/4905 DVDD:1953 X46/D0:neg 0.709092
rDVDD/4906 DVDD:1951 DVDD:1953 0.0384615
rDVDD/4907 DVDD:1951 X46/D0:neg 0.354546
rDVDD/4908 DVDD:1947 DVDD:1951 0.0384615
rDVDD/4909 DVDD:1947 DVDD:4226 0.01
rDVDD/4910 DVDD:1947 X46/D0:neg 0.709092
rDVDD/4911 DVDD:1945 DVDD:4226 0.0284615
rDVDD/4912 DVDD:1945 X46/D0:neg 0.709092
rDVDD/4913 DVDD:1943 DVDD:1945 0.0192308
rDVDD/4914 DVDD:1943 X46/D0:neg 1.04
rDVDD/4915 DVDD:1866 DVDD:4168 0.0429806
rDVDD/4916 DVDD:1859 DVDD:3994 0.119278
rDVDD/4917 DVDD:1857 DVDD:1859 0.114324
rDVDD/4918 DVDD:1855 DVDD:1857 0.114324
rDVDD/4919 DVDD:1853 DVDD:1855 0.114324
rDVDD/4920 DVDD:1851 DVDD:1853 0.114324
rDVDD/4921 DVDD:1851 DVDD:4070 0.0112703
rDVDD/4922 DVDD:1849 DVDD:4066 0.0592703
rDVDD/4923 DVDD:1849 DVDD:4052 0.0282973
rDVDD/4924 DVDD:1847 DVDD:4042 0.0422432
rDVDD/4925 DVDD:1845 DVDD:1847 0.114324
rDVDD/4926 DVDD:1843 DVDD:1845 0.114324
rDVDD/4927 DVDD:1841 DVDD:1843 0.114324
rDVDD/4928 DVDD:1839 DVDD:1841 0.114324
rDVDD/4929 DVDD:1837 DVDD:1839 0.114324
rDVDD/4930 DVDD:1835 DVDD:1837 0.114324
rDVDD/4931 DVDD:1835 DVDD:4102 0.0177568
rDVDD/4932 DVDD:1833 DVDD:4098 0.0527838
rDVDD/4933 DVDD:1833 DVDD:4084 0.0347838
rDVDD/4934 DVDD:1831 DVDD:4074 0.0357568
rDVDD/4935 DVDD:1829 DVDD:1831 0.114324
rDVDD/4936 DVDD:1827 DVDD:1829 0.114324
rDVDD/4937 DVDD:1825 DVDD:1827 0.114324
rDVDD/4938 DVDD:1823 DVDD:1825 0.114243
rDVDD/4939 DVDD:1821 DVDD:1823 0.114324
rDVDD/4940 DVDD:1819 DVDD:1821 0.114324
rDVDD/4941 DVDD:1817 DVDD:1819 0.114324
rDVDD/4942 DVDD:1817 DVDD:4134 0.0737838
rDVDD/4943 DVDD:1815 DVDD:4134 0.0405405
rDVDD/4944 DVDD:1815 DVDD:4129 1.5
rDVDD/4945 DVDD:1815 DVDD:4116 0.0908108
rDVDD/4946 DVDD:1813 DVDD:4116 0.0235135
rDVDD/4947 DVDD:1813 DVDD:4106 0.0202703
rDVDD/4948 DVDD:1811 DVDD:4106 0.0940541
rDVDD/4949 DVDD:1809 DVDD:1811 0.114324
rDVDD/4950 DVDD:1807 DVDD:1809 0.114324
rDVDD/4951 DVDD:1805 DVDD:1807 0.114324
rDVDD/4952 DVDD:1803 DVDD:1805 0.114324
rDVDD/4953 DVDD:1801 DVDD:1803 0.114324
rDVDD/4954 DVDD:1801 DVDD:4166 0.0802703
rDVDD/4955 DVDD:1799 DVDD:4166 0.0340541
rDVDD/4956 DVDD:1799 DVDD:4161 1.5
rDVDD/4957 DVDD:1799 DVDD:4148 0.0972973
rDVDD/4958 DVDD:1795 DVDD:4138 0.0875676
rDVDD/4959 DVDD:1793 DVDD:1795 0.114324
rDVDD/4960 DVDD:1791 DVDD:1793 0.114324
rDVDD/4961 DVDD:1789 DVDD:1791 0.114324
rDVDD/4962 DVDD:1787 DVDD:4182 0.0429806
rDVDD/4963 DVDD:1782 DVDD:3982 0.0252672
rDVDD/4964 DVDD:1770 DVDD:4046 0.0170426
rDVDD/4965 DVDD:1756 DVDD:4091 0.5625
rDVDD/4966 DVDD:1754 DVDD:4078 0.0132128
rDVDD/4967 DVDD:1736 DVDD:4124 0.0318351
rDVDD/4968 DVDD:1736 DVDD:4110 0.019867
rDVDD/4969 DVDD:1720 DVDD:4156 0.0280053
rDVDD/4970 DVDD:1720 DVDD:4142 0.0236968
rDVDD/4971 DVDD:1705 DVDD:3986 0.0252672
rDVDD/4972 DVDD:1693 DVDD:4048 0.0170426
rDVDD/4973 DVDD:1679 DVDD:4093 0.5625
rDVDD/4974 DVDD:1677 DVDD:4080 0.0132128
rDVDD/4975 DVDD:1659 DVDD:4126 0.0318351
rDVDD/4976 DVDD:1659 DVDD:4112 0.019867
rDVDD/4977 DVDD:1643 DVDD:4158 0.0280053
rDVDD/4978 DVDD:1643 DVDD:4144 0.0236968
rDVDD/4979 DVDD:1628 DVDD:3990 0.0252672
rDVDD/4980 DVDD:1616 DVDD:4050 0.0170426
rDVDD/4981 DVDD:1602 DVDD:4095 0.5625
rDVDD/4982 DVDD:1600 DVDD:4082 0.0132128
rDVDD/4983 DVDD:1582 DVDD:4128 0.0318351
rDVDD/4984 DVDD:1582 DVDD:4114 0.019867
rDVDD/4985 DVDD:1566 DVDD:4160 0.0280053
rDVDD/4986 DVDD:1566 DVDD:4146 0.0236968
rDVDD/4987 DVDD:1551 DVDD:3980 0.119278
rDVDD/4988 DVDD:1549 DVDD:1551 0.114324
rDVDD/4989 DVDD:1547 DVDD:1549 0.114324
rDVDD/4990 DVDD:1545 DVDD:1547 0.114324
rDVDD/4991 DVDD:1543 DVDD:1545 0.114324
rDVDD/4992 DVDD:1543 DVDD:4068 0.0112703
rDVDD/4993 DVDD:1541 DVDD:4058 0.0592703
rDVDD/4994 DVDD:1541 DVDD:4044 0.0282973
rDVDD/4995 DVDD:1539 DVDD:4040 0.0422432
rDVDD/4996 DVDD:1537 DVDD:1539 0.114324
rDVDD/4997 DVDD:1535 DVDD:1537 0.114324
rDVDD/4998 DVDD:1533 DVDD:1535 0.114324
rDVDD/4999 DVDD:1531 DVDD:1533 0.114324
rDVDD/5000 DVDD:1529 DVDD:1531 0.114324
rDVDD/5001 DVDD:1527 DVDD:1529 0.114324
rDVDD/5002 DVDD:1527 DVDD:4100 0.0177568
rDVDD/5003 DVDD:1525 DVDD:4090 0.0527838
rDVDD/5004 DVDD:1525 DVDD:4076 0.0347838
rDVDD/5005 DVDD:1523 DVDD:4072 0.0357568
rDVDD/5006 DVDD:1521 DVDD:1523 0.114324
rDVDD/5007 DVDD:1519 DVDD:1521 0.114324
rDVDD/5008 DVDD:1517 DVDD:1519 0.114324
rDVDD/5009 DVDD:1515 DVDD:1517 0.114243
rDVDD/5010 DVDD:1513 DVDD:1515 0.114324
rDVDD/5011 DVDD:1511 DVDD:1513 0.114324
rDVDD/5012 DVDD:1509 DVDD:1511 0.114324
rDVDD/5013 DVDD:1509 DVDD:4132 0.0737838
rDVDD/5014 DVDD:1507 DVDD:4132 0.0405405
rDVDD/5015 DVDD:1507 DVDD:4121 1.5
rDVDD/5016 DVDD:1507 DVDD:4108 0.0908108
rDVDD/5017 DVDD:1505 DVDD:4108 0.0235135
rDVDD/5018 DVDD:1505 DVDD:4104 0.0202703
rDVDD/5019 DVDD:1503 DVDD:4104 0.0940541
rDVDD/5020 DVDD:1501 DVDD:1503 0.114324
rDVDD/5021 DVDD:1499 DVDD:1501 0.114324
rDVDD/5022 DVDD:1497 DVDD:1499 0.114324
rDVDD/5023 DVDD:1495 DVDD:1497 0.114324
rDVDD/5024 DVDD:1493 DVDD:1495 0.114324
rDVDD/5025 DVDD:1493 DVDD:4164 0.0802703
rDVDD/5026 DVDD:1491 DVDD:4164 0.0340541
rDVDD/5027 DVDD:1491 DVDD:4153 1.5
rDVDD/5028 DVDD:1491 DVDD:4140 0.0972973
rDVDD/5029 DVDD:1487 DVDD:4136 0.0875676
rDVDD/5030 DVDD:1485 DVDD:1487 0.114324
rDVDD/5031 DVDD:1483 DVDD:1485 0.114324
rDVDD/5032 DVDD:1481 DVDD:1483 0.114324
rDVDD/5033 DVDD:1479 DVDD:1481 0.0762162
rDVDD/5034 DVDD:1479 DVDD:1866 0.0381081
rDVDD/5035 DVDD:1401 DVDD:1782 0.03375
rDVDD/5036 DVDD:1401 DVDD:1780 0.03375
rDVDD/5037 DVDD:1399 DVDD:1780 0.03375
rDVDD/5038 DVDD:1399 DVDD:1778 0.03375
rDVDD/5039 DVDD:1397 DVDD:1778 0.03375
rDVDD/5040 DVDD:1397 DVDD:1776 0.03375
rDVDD/5041 DVDD:1395 DVDD:1776 0.03375
rDVDD/5042 DVDD:1395 DVDD:1774 0.03375
rDVDD/5043 DVDD:1393 DVDD:1774 0.03375
rDVDD/5044 DVDD:1393 DVDD:4060 0.0325053
rDVDD/5045 DVDD:1391 DVDD:4060 0.0349947
rDVDD/5046 DVDD:1391 DVDD:4046 0.0167074
rDVDD/5047 DVDD:1389 DVDD:1770 0.03375
rDVDD/5048 DVDD:1389 DVDD:1768 0.03375
rDVDD/5049 DVDD:1387 DVDD:1768 0.03375
rDVDD/5050 DVDD:1387 DVDD:1766 0.03375
rDVDD/5051 DVDD:1385 DVDD:1766 0.03375
rDVDD/5052 DVDD:1385 DVDD:1764 0.03375
rDVDD/5053 DVDD:1383 DVDD:1764 0.03375
rDVDD/5054 DVDD:1383 DVDD:1762 0.03375
rDVDD/5055 DVDD:1381 DVDD:1762 0.03375
rDVDD/5056 DVDD:1381 DVDD:1760 0.03375
rDVDD/5057 DVDD:1379 DVDD:1760 0.03375
rDVDD/5058 DVDD:1379 DVDD:1758 0.03375
rDVDD/5059 DVDD:1377 DVDD:1758 0.03375
rDVDD/5060 DVDD:1377 DVDD:1756 0.03375
rDVDD/5061 DVDD:1375 DVDD:1756 0.03375
rDVDD/5062 DVDD:1375 DVDD:4078 0.0205372
rDVDD/5063 DVDD:1373 DVDD:1754 0.03375
rDVDD/5064 DVDD:1373 DVDD:1752 0.03375
rDVDD/5065 DVDD:1371 DVDD:1752 0.03375
rDVDD/5066 DVDD:1371 DVDD:1750 0.03375
rDVDD/5067 DVDD:1369 DVDD:1750 0.03375
rDVDD/5068 DVDD:1369 DVDD:1748 0.03375
rDVDD/5069 DVDD:1367 DVDD:1748 0.03375
rDVDD/5070 DVDD:1367 DVDD:1746 0.03375
rDVDD/5071 DVDD:1365 DVDD:1746 0.0337021
rDVDD/5072 DVDD:1365 DVDD:1744 0.03375
rDVDD/5073 DVDD:1363 DVDD:1744 0.03375
rDVDD/5074 DVDD:1363 DVDD:1742 0.03375
rDVDD/5075 DVDD:1361 DVDD:1742 0.03375
rDVDD/5076 DVDD:1361 DVDD:1740 0.03375
rDVDD/5077 DVDD:1359 DVDD:1740 0.03375
rDVDD/5078 DVDD:1359 DVDD:1738 0.03375
rDVDD/5079 DVDD:1357 DVDD:1738 0.03375
rDVDD/5080 DVDD:1357 DVDD:4124 0.00191489
rDVDD/5081 DVDD:1355 DVDD:4110 0.013883
rDVDD/5082 DVDD:1355 DVDD:1734 0.03375
rDVDD/5083 DVDD:1353 DVDD:1734 0.03375
rDVDD/5084 DVDD:1353 DVDD:1732 0.03375
rDVDD/5085 DVDD:1351 DVDD:1732 0.03375
rDVDD/5086 DVDD:1351 DVDD:1730 0.03375
rDVDD/5087 DVDD:1349 DVDD:1730 0.03375
rDVDD/5088 DVDD:1349 DVDD:1728 0.03375
rDVDD/5089 DVDD:1347 DVDD:1728 0.03375
rDVDD/5090 DVDD:1347 DVDD:1726 0.03375
rDVDD/5091 DVDD:1345 DVDD:1726 0.03375
rDVDD/5092 DVDD:1345 DVDD:1724 0.03375
rDVDD/5093 DVDD:1343 DVDD:1724 0.03375
rDVDD/5094 DVDD:1343 DVDD:1722 0.03375
rDVDD/5095 DVDD:1341 DVDD:1722 0.03375
rDVDD/5096 DVDD:1341 DVDD:4156 0.00574468
rDVDD/5097 DVDD:1339 DVDD:4142 0.0100532
rDVDD/5098 DVDD:1339 DVDD:1718 0.03375
rDVDD/5099 DVDD:1337 DVDD:1718 0.03375
rDVDD/5100 DVDD:1337 DVDD:1716 0.03375
rDVDD/5101 DVDD:1335 DVDD:1716 0.03375
rDVDD/5102 DVDD:1335 DVDD:1714 0.03375
rDVDD/5103 DVDD:1333 DVDD:1714 0.03375
rDVDD/5104 DVDD:1333 DVDD:1712 0.03375
rDVDD/5105 DVDD:1331 DVDD:1712 0.03375
rDVDD/5106 DVDD:1331 DVDD:1710 0.03375
rDVDD/5107 DVDD:1329 DVDD:1710 0.01125
rDVDD/5108 DVDD:1329 DVDD:4170 0.0364693
rDVDD/5109 DVDD:1251 DVDD:1705 0.03375
rDVDD/5110 DVDD:1251 DVDD:1703 0.03375
rDVDD/5111 DVDD:1249 DVDD:1703 0.03375
rDVDD/5112 DVDD:1249 DVDD:1701 0.03375
rDVDD/5113 DVDD:1247 DVDD:1701 0.03375
rDVDD/5114 DVDD:1247 DVDD:1699 0.03375
rDVDD/5115 DVDD:1245 DVDD:1699 0.03375
rDVDD/5116 DVDD:1245 DVDD:1697 0.03375
rDVDD/5117 DVDD:1243 DVDD:1697 0.03375
rDVDD/5118 DVDD:1243 DVDD:4062 0.0325053
rDVDD/5119 DVDD:1241 DVDD:4062 0.0349947
rDVDD/5120 DVDD:1241 DVDD:4048 0.0167074
rDVDD/5121 DVDD:1239 DVDD:1693 0.03375
rDVDD/5122 DVDD:1239 DVDD:1691 0.03375
rDVDD/5123 DVDD:1237 DVDD:1691 0.03375
rDVDD/5124 DVDD:1237 DVDD:1689 0.03375
rDVDD/5125 DVDD:1235 DVDD:1689 0.03375
rDVDD/5126 DVDD:1235 DVDD:1687 0.03375
rDVDD/5127 DVDD:1233 DVDD:1687 0.03375
rDVDD/5128 DVDD:1233 DVDD:1685 0.03375
rDVDD/5129 DVDD:1231 DVDD:1685 0.03375
rDVDD/5130 DVDD:1231 DVDD:1683 0.03375
rDVDD/5131 DVDD:1229 DVDD:1683 0.03375
rDVDD/5132 DVDD:1229 DVDD:1681 0.03375
rDVDD/5133 DVDD:1227 DVDD:1681 0.03375
rDVDD/5134 DVDD:1227 DVDD:1679 0.03375
rDVDD/5135 DVDD:1225 DVDD:1679 0.03375
rDVDD/5136 DVDD:1225 DVDD:4080 0.0205372
rDVDD/5137 DVDD:1223 DVDD:1677 0.03375
rDVDD/5138 DVDD:1223 DVDD:1675 0.03375
rDVDD/5139 DVDD:1221 DVDD:1675 0.03375
rDVDD/5140 DVDD:1221 DVDD:1673 0.03375
rDVDD/5141 DVDD:1219 DVDD:1673 0.03375
rDVDD/5142 DVDD:1219 DVDD:1671 0.03375
rDVDD/5143 DVDD:1217 DVDD:1671 0.03375
rDVDD/5144 DVDD:1217 DVDD:1669 0.03375
rDVDD/5145 DVDD:1215 DVDD:1669 0.0337021
rDVDD/5146 DVDD:1215 DVDD:1667 0.03375
rDVDD/5147 DVDD:1213 DVDD:1667 0.03375
rDVDD/5148 DVDD:1213 DVDD:1665 0.03375
rDVDD/5149 DVDD:1211 DVDD:1665 0.03375
rDVDD/5150 DVDD:1211 DVDD:1663 0.03375
rDVDD/5151 DVDD:1209 DVDD:1663 0.03375
rDVDD/5152 DVDD:1209 DVDD:1661 0.03375
rDVDD/5153 DVDD:1207 DVDD:1661 0.03375
rDVDD/5154 DVDD:1207 DVDD:4126 0.00191489
rDVDD/5155 DVDD:1205 DVDD:4112 0.013883
rDVDD/5156 DVDD:1205 DVDD:1657 0.03375
rDVDD/5157 DVDD:1203 DVDD:1657 0.03375
rDVDD/5158 DVDD:1203 DVDD:1655 0.03375
rDVDD/5159 DVDD:1201 DVDD:1655 0.03375
rDVDD/5160 DVDD:1201 DVDD:1653 0.03375
rDVDD/5161 DVDD:1199 DVDD:1653 0.03375
rDVDD/5162 DVDD:1199 DVDD:1651 0.03375
rDVDD/5163 DVDD:1197 DVDD:1651 0.03375
rDVDD/5164 DVDD:1197 DVDD:1649 0.03375
rDVDD/5165 DVDD:1195 DVDD:1649 0.03375
rDVDD/5166 DVDD:1195 DVDD:1647 0.03375
rDVDD/5167 DVDD:1193 DVDD:1647 0.03375
rDVDD/5168 DVDD:1193 DVDD:1645 0.03375
rDVDD/5169 DVDD:1191 DVDD:1645 0.03375
rDVDD/5170 DVDD:1191 DVDD:4158 0.00574468
rDVDD/5171 DVDD:1189 DVDD:4144 0.0100532
rDVDD/5172 DVDD:1189 DVDD:1641 0.03375
rDVDD/5173 DVDD:1187 DVDD:1641 0.03375
rDVDD/5174 DVDD:1187 DVDD:1639 0.03375
rDVDD/5175 DVDD:1185 DVDD:1639 0.03375
rDVDD/5176 DVDD:1185 DVDD:1637 0.03375
rDVDD/5177 DVDD:1183 DVDD:1637 0.03375
rDVDD/5178 DVDD:1183 DVDD:1635 0.03375
rDVDD/5179 DVDD:1181 DVDD:1635 0.03375
rDVDD/5180 DVDD:1181 DVDD:1633 0.03375
rDVDD/5181 DVDD:1179 DVDD:1633 0.01125
rDVDD/5182 DVDD:1179 DVDD:4174 0.0364693
rDVDD/5183 DVDD:1101 DVDD:1628 0.03375
rDVDD/5184 DVDD:1101 DVDD:1626 0.03375
rDVDD/5185 DVDD:1099 DVDD:1626 0.03375
rDVDD/5186 DVDD:1099 DVDD:1624 0.03375
rDVDD/5187 DVDD:1097 DVDD:1624 0.03375
rDVDD/5188 DVDD:1097 DVDD:1622 0.03375
rDVDD/5189 DVDD:1095 DVDD:1622 0.03375
rDVDD/5190 DVDD:1095 DVDD:1620 0.03375
rDVDD/5191 DVDD:1093 DVDD:1620 0.03375
rDVDD/5192 DVDD:1093 DVDD:4064 0.0325053
rDVDD/5193 DVDD:1091 DVDD:4064 0.0349947
rDVDD/5194 DVDD:1091 DVDD:4050 0.0167074
rDVDD/5195 DVDD:1089 DVDD:1616 0.03375
rDVDD/5196 DVDD:1089 DVDD:1614 0.03375
rDVDD/5197 DVDD:1087 DVDD:1614 0.03375
rDVDD/5198 DVDD:1087 DVDD:1612 0.03375
rDVDD/5199 DVDD:1085 DVDD:1612 0.03375
rDVDD/5200 DVDD:1085 DVDD:1610 0.03375
rDVDD/5201 DVDD:1083 DVDD:1610 0.03375
rDVDD/5202 DVDD:1083 DVDD:1608 0.03375
rDVDD/5203 DVDD:1081 DVDD:1608 0.03375
rDVDD/5204 DVDD:1081 DVDD:1606 0.03375
rDVDD/5205 DVDD:1079 DVDD:1606 0.03375
rDVDD/5206 DVDD:1079 DVDD:1604 0.03375
rDVDD/5207 DVDD:1077 DVDD:1604 0.03375
rDVDD/5208 DVDD:1077 DVDD:1602 0.03375
rDVDD/5209 DVDD:1075 DVDD:1602 0.03375
rDVDD/5210 DVDD:1075 DVDD:4082 0.0205372
rDVDD/5211 DVDD:1073 DVDD:1600 0.03375
rDVDD/5212 DVDD:1073 DVDD:1598 0.03375
rDVDD/5213 DVDD:1071 DVDD:1598 0.03375
rDVDD/5214 DVDD:1071 DVDD:1596 0.03375
rDVDD/5215 DVDD:1069 DVDD:1596 0.03375
rDVDD/5216 DVDD:1069 DVDD:1594 0.03375
rDVDD/5217 DVDD:1067 DVDD:1594 0.03375
rDVDD/5218 DVDD:1067 DVDD:1592 0.03375
rDVDD/5219 DVDD:1065 DVDD:1592 0.0337021
rDVDD/5220 DVDD:1065 DVDD:1590 0.03375
rDVDD/5221 DVDD:1063 DVDD:1590 0.03375
rDVDD/5222 DVDD:1063 DVDD:1588 0.03375
rDVDD/5223 DVDD:1061 DVDD:1588 0.03375
rDVDD/5224 DVDD:1061 DVDD:1586 0.03375
rDVDD/5225 DVDD:1059 DVDD:1586 0.03375
rDVDD/5226 DVDD:1059 DVDD:1584 0.03375
rDVDD/5227 DVDD:1057 DVDD:1584 0.03375
rDVDD/5228 DVDD:1057 DVDD:4128 0.00191489
rDVDD/5229 DVDD:1055 DVDD:4114 0.013883
rDVDD/5230 DVDD:1055 DVDD:1580 0.03375
rDVDD/5231 DVDD:1053 DVDD:1580 0.03375
rDVDD/5232 DVDD:1053 DVDD:1578 0.03375
rDVDD/5233 DVDD:1051 DVDD:1578 0.03375
rDVDD/5234 DVDD:1051 DVDD:1576 0.03375
rDVDD/5235 DVDD:1049 DVDD:1576 0.03375
rDVDD/5236 DVDD:1049 DVDD:1574 0.03375
rDVDD/5237 DVDD:1047 DVDD:1574 0.03375
rDVDD/5238 DVDD:1047 DVDD:1572 0.03375
rDVDD/5239 DVDD:1045 DVDD:1572 0.03375
rDVDD/5240 DVDD:1045 DVDD:1570 0.03375
rDVDD/5241 DVDD:1043 DVDD:1570 0.03375
rDVDD/5242 DVDD:1043 DVDD:1568 0.03375
rDVDD/5243 DVDD:1041 DVDD:1568 0.03375
rDVDD/5244 DVDD:1041 DVDD:4160 0.00574468
rDVDD/5245 DVDD:1039 DVDD:4146 0.0100532
rDVDD/5246 DVDD:1039 DVDD:1564 0.03375
rDVDD/5247 DVDD:1037 DVDD:1564 0.03375
rDVDD/5248 DVDD:1037 DVDD:1562 0.03375
rDVDD/5249 DVDD:1035 DVDD:1562 0.03375
rDVDD/5250 DVDD:1035 DVDD:1560 0.03375
rDVDD/5251 DVDD:1033 DVDD:1560 0.03375
rDVDD/5252 DVDD:1033 DVDD:1558 0.03375
rDVDD/5253 DVDD:1031 DVDD:1558 0.03375
rDVDD/5254 DVDD:1031 DVDD:1556 0.03375
rDVDD/5255 DVDD:1029 DVDD:1556 0.01125
rDVDD/5256 DVDD:1029 DVDD:4178 0.0364693
rDVDD/5257 DVDD:954 DVDD:1789 0.0762162
rDVDD/5258 DVDD:954 DVDD:1787 0.0381081
rDVDD/5259 X46/X30/D0:neg DVDD:4202 1.73333
rDVDD/5260 X46/X30/D0:neg DVDD:4192 1.73333
rDVDD/5261 X46/X30/D0:neg DVDD:4182 5.2
rDVDD/5262 X46/X30/D0:neg DVDD:4178 1.3
rDVDD/5263 X46/X30/D0:neg DVDD:4174 1.3
rDVDD/5264 X46/X30/D0:neg DVDD:4170 1.3
rDVDD/5265 X46/X30/D0:neg DVDD:4168 5.2
rDVDD/5266 X46/X30/D0:neg DVDD:4148 0.866667
rDVDD/5267 X46/X30/D0:neg DVDD:4140 0.866667
rDVDD/5268 X46/X30/D0:neg DVDD:4064 1.73333
rDVDD/5269 X46/X30/D0:neg DVDD:4062 1.73333
rDVDD/5270 X46/X30/D0:neg DVDD:4060 1.73333
rDVDD/5271 X46/X30/D0:neg DVDD:4034 1.73333
rDVDD/5272 X46/X30/D0:neg DVDD:4024 1.73333
rDVDD/5273 X46/X30/D0:neg DVDD:3994 1.73333
rDVDD/5274 X46/X30/D0:neg DVDD:3990 1.73333
rDVDD/5275 X46/X30/D0:neg DVDD:3986 1.73333
rDVDD/5276 X46/X30/D0:neg DVDD:3982 1.73333
rDVDD/5277 X46/X30/D0:neg DVDD:3980 1.73333
rDVDD/5278 X46/X30/D0:neg DVDD:1866 1.73333
rDVDD/5279 X46/X30/D0:neg DVDD:1859 0.866667
rDVDD/5280 X46/X30/D0:neg DVDD:1857 0.866667
rDVDD/5281 X46/X30/D0:neg DVDD:1855 0.866667
rDVDD/5282 X46/X30/D0:neg DVDD:1853 0.866667
rDVDD/5283 X46/X30/D0:neg DVDD:1851 0.866667
rDVDD/5284 X46/X30/D0:neg DVDD:1849 0.866667
rDVDD/5285 X46/X30/D0:neg DVDD:1847 0.866667
rDVDD/5286 X46/X30/D0:neg DVDD:1845 0.866667
rDVDD/5287 X46/X30/D0:neg DVDD:1843 0.866667
rDVDD/5288 X46/X30/D0:neg DVDD:1841 0.866667
rDVDD/5289 X46/X30/D0:neg DVDD:1839 0.866667
rDVDD/5290 X46/X30/D0:neg DVDD:1837 0.866667
rDVDD/5291 X46/X30/D0:neg DVDD:1835 0.866667
rDVDD/5292 X46/X30/D0:neg DVDD:1833 0.866667
rDVDD/5293 X46/X30/D0:neg DVDD:1831 0.866667
rDVDD/5294 X46/X30/D0:neg DVDD:1829 0.866667
rDVDD/5295 X46/X30/D0:neg DVDD:1827 0.866667
rDVDD/5296 X46/X30/D0:neg DVDD:1825 0.866667
rDVDD/5297 X46/X30/D0:neg DVDD:1823 0.866667
rDVDD/5298 X46/X30/D0:neg DVDD:1821 0.866667
rDVDD/5299 X46/X30/D0:neg DVDD:1819 0.866667
rDVDD/5300 X46/X30/D0:neg DVDD:1817 0.866667
rDVDD/5301 X46/X30/D0:neg DVDD:1815 0.866667
rDVDD/5302 X46/X30/D0:neg DVDD:1813 0.866667
rDVDD/5303 X46/X30/D0:neg DVDD:1811 0.866667
rDVDD/5304 X46/X30/D0:neg DVDD:1809 0.866667
rDVDD/5305 X46/X30/D0:neg DVDD:1807 0.866667
rDVDD/5306 X46/X30/D0:neg DVDD:1805 0.866667
rDVDD/5307 X46/X30/D0:neg DVDD:1803 0.866667
rDVDD/5308 X46/X30/D0:neg DVDD:1801 0.866667
rDVDD/5309 X46/X30/D0:neg DVDD:1799 0.866667
rDVDD/5310 X46/X30/D0:neg DVDD:1795 0.866667
rDVDD/5311 X46/X30/D0:neg DVDD:1793 0.866667
rDVDD/5312 X46/X30/D0:neg DVDD:1791 0.866667
rDVDD/5313 X46/X30/D0:neg DVDD:1789 0.866667
rDVDD/5314 X46/X30/D0:neg DVDD:1787 1.73333
rDVDD/5315 X46/X30/D0:neg DVDD:1782 1.73333
rDVDD/5316 X46/X30/D0:neg DVDD:1780 1.73333
rDVDD/5317 X46/X30/D0:neg DVDD:1778 1.73333
rDVDD/5318 X46/X30/D0:neg DVDD:1776 1.73333
rDVDD/5319 X46/X30/D0:neg DVDD:1774 1.73333
rDVDD/5320 X46/X30/D0:neg DVDD:1770 1.73333
rDVDD/5321 X46/X30/D0:neg DVDD:1768 1.73333
rDVDD/5322 X46/X30/D0:neg DVDD:1766 1.73333
rDVDD/5323 X46/X30/D0:neg DVDD:1764 1.73333
rDVDD/5324 X46/X30/D0:neg DVDD:1762 1.73333
rDVDD/5325 X46/X30/D0:neg DVDD:1760 1.73333
rDVDD/5326 X46/X30/D0:neg DVDD:1758 1.73333
rDVDD/5327 X46/X30/D0:neg DVDD:1756 1.73333
rDVDD/5328 X46/X30/D0:neg DVDD:1754 1.73333
rDVDD/5329 X46/X30/D0:neg DVDD:1752 1.73333
rDVDD/5330 X46/X30/D0:neg DVDD:1750 1.73333
rDVDD/5331 X46/X30/D0:neg DVDD:1748 1.73333
rDVDD/5332 X46/X30/D0:neg DVDD:1746 1.73333
rDVDD/5333 X46/X30/D0:neg DVDD:1744 1.73333
rDVDD/5334 X46/X30/D0:neg DVDD:1742 1.73333
rDVDD/5335 X46/X30/D0:neg DVDD:1740 1.73333
rDVDD/5336 X46/X30/D0:neg DVDD:1738 1.73333
rDVDD/5337 X46/X30/D0:neg DVDD:1736 1.73333
rDVDD/5338 X46/X30/D0:neg DVDD:1734 1.73333
rDVDD/5339 X46/X30/D0:neg DVDD:1732 1.73333
rDVDD/5340 X46/X30/D0:neg DVDD:1730 1.73333
rDVDD/5341 X46/X30/D0:neg DVDD:1728 1.73333
rDVDD/5342 X46/X30/D0:neg DVDD:1726 1.73333
rDVDD/5343 X46/X30/D0:neg DVDD:1724 1.73333
rDVDD/5344 X46/X30/D0:neg DVDD:1722 1.73333
rDVDD/5345 X46/X30/D0:neg DVDD:1720 1.73333
rDVDD/5346 X46/X30/D0:neg DVDD:1718 1.73333
rDVDD/5347 X46/X30/D0:neg DVDD:1716 1.73333
rDVDD/5348 X46/X30/D0:neg DVDD:1714 1.73333
rDVDD/5349 X46/X30/D0:neg DVDD:1712 1.73333
rDVDD/5350 X46/X30/D0:neg DVDD:1710 1.73333
rDVDD/5351 X46/X30/D0:neg DVDD:1705 1.73333
rDVDD/5352 X46/X30/D0:neg DVDD:1703 1.73333
rDVDD/5353 X46/X30/D0:neg DVDD:1701 1.73333
rDVDD/5354 X46/X30/D0:neg DVDD:1699 1.73333
rDVDD/5355 X46/X30/D0:neg DVDD:1697 1.73333
rDVDD/5356 X46/X30/D0:neg DVDD:1693 1.73333
rDVDD/5357 X46/X30/D0:neg DVDD:1691 1.73333
rDVDD/5358 X46/X30/D0:neg DVDD:1689 1.73333
rDVDD/5359 X46/X30/D0:neg DVDD:1687 1.73333
rDVDD/5360 X46/X30/D0:neg DVDD:1685 1.73333
rDVDD/5361 X46/X30/D0:neg DVDD:1683 1.73333
rDVDD/5362 X46/X30/D0:neg DVDD:1681 1.73333
rDVDD/5363 X46/X30/D0:neg DVDD:1679 1.73333
rDVDD/5364 X46/X30/D0:neg DVDD:1677 1.73333
rDVDD/5365 X46/X30/D0:neg DVDD:1675 1.73333
rDVDD/5366 X46/X30/D0:neg DVDD:1673 1.73333
rDVDD/5367 X46/X30/D0:neg DVDD:1671 1.73333
rDVDD/5368 X46/X30/D0:neg DVDD:1669 1.73333
rDVDD/5369 X46/X30/D0:neg DVDD:1667 1.73333
rDVDD/5370 X46/X30/D0:neg DVDD:1665 1.73333
rDVDD/5371 X46/X30/D0:neg DVDD:1663 1.73333
rDVDD/5372 X46/X30/D0:neg DVDD:1661 1.73333
rDVDD/5373 X46/X30/D0:neg DVDD:1659 1.73333
rDVDD/5374 X46/X30/D0:neg DVDD:1657 1.73333
rDVDD/5375 X46/X30/D0:neg DVDD:1655 1.73333
rDVDD/5376 X46/X30/D0:neg DVDD:1653 1.73333
rDVDD/5377 X46/X30/D0:neg DVDD:1651 1.73333
rDVDD/5378 X46/X30/D0:neg DVDD:1649 1.73333
rDVDD/5379 X46/X30/D0:neg DVDD:1647 1.73333
rDVDD/5380 X46/X30/D0:neg DVDD:1645 1.73333
rDVDD/5381 X46/X30/D0:neg DVDD:1643 1.73333
rDVDD/5382 X46/X30/D0:neg DVDD:1641 1.73333
rDVDD/5383 X46/X30/D0:neg DVDD:1639 1.73333
rDVDD/5384 X46/X30/D0:neg DVDD:1637 1.73333
rDVDD/5385 X46/X30/D0:neg DVDD:1635 1.73333
rDVDD/5386 X46/X30/D0:neg DVDD:1633 1.73333
rDVDD/5387 X46/X30/D0:neg DVDD:1628 1.73333
rDVDD/5388 X46/X30/D0:neg DVDD:1626 1.73333
rDVDD/5389 X46/X30/D0:neg DVDD:1624 1.73333
rDVDD/5390 X46/X30/D0:neg DVDD:1622 1.73333
rDVDD/5391 X46/X30/D0:neg DVDD:1620 1.73333
rDVDD/5392 X46/X30/D0:neg DVDD:1616 1.73333
rDVDD/5393 X46/X30/D0:neg DVDD:1614 1.73333
rDVDD/5394 X46/X30/D0:neg DVDD:1612 1.73333
rDVDD/5395 X46/X30/D0:neg DVDD:1610 1.73333
rDVDD/5396 X46/X30/D0:neg DVDD:1608 1.73333
rDVDD/5397 X46/X30/D0:neg DVDD:1606 1.73333
rDVDD/5398 X46/X30/D0:neg DVDD:1604 1.73333
rDVDD/5399 X46/X30/D0:neg DVDD:1602 1.73333
rDVDD/5400 X46/X30/D0:neg DVDD:1600 1.73333
rDVDD/5401 X46/X30/D0:neg DVDD:1598 1.73333
rDVDD/5402 X46/X30/D0:neg DVDD:1596 1.73333
rDVDD/5403 X46/X30/D0:neg DVDD:1594 1.73333
rDVDD/5404 X46/X30/D0:neg DVDD:1592 1.73333
rDVDD/5405 X46/X30/D0:neg DVDD:1590 1.73333
rDVDD/5406 X46/X30/D0:neg DVDD:1588 1.73333
rDVDD/5407 X46/X30/D0:neg DVDD:1586 1.73333
rDVDD/5408 X46/X30/D0:neg DVDD:1584 1.73333
rDVDD/5409 X46/X30/D0:neg DVDD:1582 1.73333
rDVDD/5410 X46/X30/D0:neg DVDD:1580 1.73333
rDVDD/5411 X46/X30/D0:neg DVDD:1578 1.73333
rDVDD/5412 X46/X30/D0:neg DVDD:1576 1.73333
rDVDD/5413 X46/X30/D0:neg DVDD:1574 1.73333
rDVDD/5414 X46/X30/D0:neg DVDD:1572 1.73333
rDVDD/5415 X46/X30/D0:neg DVDD:1570 1.73333
rDVDD/5416 X46/X30/D0:neg DVDD:1568 1.73333
rDVDD/5417 X46/X30/D0:neg DVDD:1566 1.73333
rDVDD/5418 X46/X30/D0:neg DVDD:1564 1.73333
rDVDD/5419 X46/X30/D0:neg DVDD:1562 1.73333
rDVDD/5420 X46/X30/D0:neg DVDD:1560 1.73333
rDVDD/5421 X46/X30/D0:neg DVDD:1558 1.73333
rDVDD/5422 X46/X30/D0:neg DVDD:1556 1.73333
rDVDD/5423 X46/X30/D0:neg DVDD:1551 0.866667
rDVDD/5424 X46/X30/D0:neg DVDD:1549 0.866667
rDVDD/5425 X46/X30/D0:neg DVDD:1547 0.866667
rDVDD/5426 X46/X30/D0:neg DVDD:1545 0.866667
rDVDD/5427 X46/X30/D0:neg DVDD:1543 0.866667
rDVDD/5428 X46/X30/D0:neg DVDD:1541 0.866667
rDVDD/5429 X46/X30/D0:neg DVDD:1539 0.866667
rDVDD/5430 X46/X30/D0:neg DVDD:1537 0.866667
rDVDD/5431 X46/X30/D0:neg DVDD:1535 0.866667
rDVDD/5432 X46/X30/D0:neg DVDD:1533 0.866667
rDVDD/5433 X46/X30/D0:neg DVDD:1531 0.866667
rDVDD/5434 X46/X30/D0:neg DVDD:1529 0.866667
rDVDD/5435 X46/X30/D0:neg DVDD:1527 0.866667
rDVDD/5436 X46/X30/D0:neg DVDD:1525 0.866667
rDVDD/5437 X46/X30/D0:neg DVDD:1523 0.866667
rDVDD/5438 X46/X30/D0:neg DVDD:1521 0.866667
rDVDD/5439 X46/X30/D0:neg DVDD:1519 0.866667
rDVDD/5440 X46/X30/D0:neg DVDD:1517 0.866667
rDVDD/5441 X46/X30/D0:neg DVDD:1515 0.866667
rDVDD/5442 X46/X30/D0:neg DVDD:1513 0.866667
rDVDD/5443 X46/X30/D0:neg DVDD:1511 0.866667
rDVDD/5444 X46/X30/D0:neg DVDD:1509 0.866667
rDVDD/5445 X46/X30/D0:neg DVDD:1507 0.866667
rDVDD/5446 X46/X30/D0:neg DVDD:1505 0.866667
rDVDD/5447 X46/X30/D0:neg DVDD:1503 0.866667
rDVDD/5448 X46/X30/D0:neg DVDD:1501 0.866667
rDVDD/5449 X46/X30/D0:neg DVDD:1499 0.866667
rDVDD/5450 X46/X30/D0:neg DVDD:1497 0.866667
rDVDD/5451 X46/X30/D0:neg DVDD:1495 0.866667
rDVDD/5452 X46/X30/D0:neg DVDD:1493 0.866667
rDVDD/5453 X46/X30/D0:neg DVDD:1491 0.866667
rDVDD/5454 X46/X30/D0:neg DVDD:1487 0.866667
rDVDD/5455 X46/X30/D0:neg DVDD:1485 0.866667
rDVDD/5456 X46/X30/D0:neg DVDD:1483 0.866667
rDVDD/5457 X46/X30/D0:neg DVDD:1481 0.866667
rDVDD/5458 X46/X30/D0:neg DVDD:1479 5.2
rDVDD/5459 X46/X30/D0:neg DVDD:1401 0.866667
rDVDD/5460 X46/X30/D0:neg DVDD:1399 0.866667
rDVDD/5461 X46/X30/D0:neg DVDD:1397 0.866667
rDVDD/5462 X46/X30/D0:neg DVDD:1395 0.866667
rDVDD/5463 X46/X30/D0:neg DVDD:1393 0.866667
rDVDD/5464 X46/X30/D0:neg DVDD:1391 0.866667
rDVDD/5465 X46/X30/D0:neg DVDD:1389 0.866667
rDVDD/5466 X46/X30/D0:neg DVDD:1387 0.866667
rDVDD/5467 X46/X30/D0:neg DVDD:1385 0.866667
rDVDD/5468 X46/X30/D0:neg DVDD:1383 0.866667
rDVDD/5469 X46/X30/D0:neg DVDD:1381 0.866667
rDVDD/5470 X46/X30/D0:neg DVDD:1379 0.866667
rDVDD/5471 X46/X30/D0:neg DVDD:1377 0.866667
rDVDD/5472 X46/X30/D0:neg DVDD:1375 0.866667
rDVDD/5473 X46/X30/D0:neg DVDD:1373 0.866667
rDVDD/5474 X46/X30/D0:neg DVDD:1371 0.866667
rDVDD/5475 X46/X30/D0:neg DVDD:1369 0.866667
rDVDD/5476 X46/X30/D0:neg DVDD:1367 0.866667
rDVDD/5477 X46/X30/D0:neg DVDD:1365 0.866667
rDVDD/5478 X46/X30/D0:neg DVDD:1363 0.866667
rDVDD/5479 X46/X30/D0:neg DVDD:1361 0.866667
rDVDD/5480 X46/X30/D0:neg DVDD:1359 0.866667
rDVDD/5481 X46/X30/D0:neg DVDD:1357 0.866667
rDVDD/5482 X46/X30/D0:neg DVDD:1355 0.866667
rDVDD/5483 X46/X30/D0:neg DVDD:1353 0.866667
rDVDD/5484 X46/X30/D0:neg DVDD:1351 0.866667
rDVDD/5485 X46/X30/D0:neg DVDD:1349 0.866667
rDVDD/5486 X46/X30/D0:neg DVDD:1347 0.866667
rDVDD/5487 X46/X30/D0:neg DVDD:1345 0.866667
rDVDD/5488 X46/X30/D0:neg DVDD:1343 0.866667
rDVDD/5489 X46/X30/D0:neg DVDD:1341 0.866667
rDVDD/5490 X46/X30/D0:neg DVDD:1339 0.866667
rDVDD/5491 X46/X30/D0:neg DVDD:1337 0.866667
rDVDD/5492 X46/X30/D0:neg DVDD:1335 0.866667
rDVDD/5493 X46/X30/D0:neg DVDD:1333 0.866667
rDVDD/5494 X46/X30/D0:neg DVDD:1331 0.866667
rDVDD/5495 X46/X30/D0:neg DVDD:1329 2.6
rDVDD/5496 X46/X30/D0:neg DVDD:1251 0.866667
rDVDD/5497 X46/X30/D0:neg DVDD:1249 0.866667
rDVDD/5498 X46/X30/D0:neg DVDD:1247 0.866667
rDVDD/5499 X46/X30/D0:neg DVDD:1245 0.866667
rDVDD/5500 X46/X30/D0:neg DVDD:1243 0.866667
rDVDD/5501 X46/X30/D0:neg DVDD:1241 0.866667
rDVDD/5502 X46/X30/D0:neg DVDD:1239 0.866667
rDVDD/5503 X46/X30/D0:neg DVDD:1237 0.866667
rDVDD/5504 X46/X30/D0:neg DVDD:1235 0.866667
rDVDD/5505 X46/X30/D0:neg DVDD:1233 0.866667
rDVDD/5506 X46/X30/D0:neg DVDD:1231 0.866667
rDVDD/5507 X46/X30/D0:neg DVDD:1229 0.866667
rDVDD/5508 X46/X30/D0:neg DVDD:1227 0.866667
rDVDD/5509 X46/X30/D0:neg DVDD:1225 0.866667
rDVDD/5510 X46/X30/D0:neg DVDD:1223 0.866667
rDVDD/5511 X46/X30/D0:neg DVDD:1221 0.866667
rDVDD/5512 X46/X30/D0:neg DVDD:1219 0.866667
rDVDD/5513 X46/X30/D0:neg DVDD:1217 0.866667
rDVDD/5514 X46/X30/D0:neg DVDD:1215 0.866667
rDVDD/5515 X46/X30/D0:neg DVDD:1213 0.866667
rDVDD/5516 X46/X30/D0:neg DVDD:1211 0.866667
rDVDD/5517 X46/X30/D0:neg DVDD:1209 0.866667
rDVDD/5518 X46/X30/D0:neg DVDD:1207 0.866667
rDVDD/5519 X46/X30/D0:neg DVDD:1205 0.866667
rDVDD/5520 X46/X30/D0:neg DVDD:1203 0.866667
rDVDD/5521 X46/X30/D0:neg DVDD:1201 0.866667
rDVDD/5522 X46/X30/D0:neg DVDD:1199 0.866667
rDVDD/5523 X46/X30/D0:neg DVDD:1197 0.866667
rDVDD/5524 X46/X30/D0:neg DVDD:1195 0.866667
rDVDD/5525 X46/X30/D0:neg DVDD:1193 0.866667
rDVDD/5526 X46/X30/D0:neg DVDD:1191 0.866667
rDVDD/5527 X46/X30/D0:neg DVDD:1189 0.866667
rDVDD/5528 X46/X30/D0:neg DVDD:1187 0.866667
rDVDD/5529 X46/X30/D0:neg DVDD:1185 0.866667
rDVDD/5530 X46/X30/D0:neg DVDD:1183 0.866667
rDVDD/5531 X46/X30/D0:neg DVDD:1181 0.866667
rDVDD/5532 X46/X30/D0:neg DVDD:1179 2.6
rDVDD/5533 X46/X30/D0:neg DVDD:1101 0.866667
rDVDD/5534 X46/X30/D0:neg DVDD:1099 0.866667
rDVDD/5535 X46/X30/D0:neg DVDD:1097 0.866667
rDVDD/5536 X46/X30/D0:neg DVDD:1095 0.866667
rDVDD/5537 X46/X30/D0:neg DVDD:1093 0.866667
rDVDD/5538 X46/X30/D0:neg DVDD:1091 0.866667
rDVDD/5539 X46/X30/D0:neg DVDD:1089 0.866667
rDVDD/5540 X46/X30/D0:neg DVDD:1087 0.866667
rDVDD/5541 X46/X30/D0:neg DVDD:1085 0.866667
rDVDD/5542 X46/X30/D0:neg DVDD:1083 0.866667
rDVDD/5543 X46/X30/D0:neg DVDD:1081 0.866667
rDVDD/5544 X46/X30/D0:neg DVDD:1079 0.866667
rDVDD/5545 X46/X30/D0:neg DVDD:1077 0.866667
rDVDD/5546 X46/X30/D0:neg DVDD:1075 0.866667
rDVDD/5547 X46/X30/D0:neg DVDD:1073 0.866667
rDVDD/5548 X46/X30/D0:neg DVDD:1071 0.866667
rDVDD/5549 X46/X30/D0:neg DVDD:1069 0.866667
rDVDD/5550 X46/X30/D0:neg DVDD:1067 0.866667
rDVDD/5551 X46/X30/D0:neg DVDD:1065 0.866667
rDVDD/5552 X46/X30/D0:neg DVDD:1063 0.866667
rDVDD/5553 X46/X30/D0:neg DVDD:1061 0.866667
rDVDD/5554 X46/X30/D0:neg DVDD:1059 0.866667
rDVDD/5555 X46/X30/D0:neg DVDD:1057 0.866667
rDVDD/5556 X46/X30/D0:neg DVDD:1055 0.866667
rDVDD/5557 X46/X30/D0:neg DVDD:1053 0.866667
rDVDD/5558 X46/X30/D0:neg DVDD:1051 0.866667
rDVDD/5559 X46/X30/D0:neg DVDD:1049 0.866667
rDVDD/5560 X46/X30/D0:neg DVDD:1047 0.866667
rDVDD/5561 X46/X30/D0:neg DVDD:1045 0.866667
rDVDD/5562 X46/X30/D0:neg DVDD:1043 0.866667
rDVDD/5563 X46/X30/D0:neg DVDD:1041 0.866667
rDVDD/5564 X46/X30/D0:neg DVDD:1039 0.866667
rDVDD/5565 X46/X30/D0:neg DVDD:1037 0.866667
rDVDD/5566 X46/X30/D0:neg DVDD:1035 0.866667
rDVDD/5567 X46/X30/D0:neg DVDD:1033 0.866667
rDVDD/5568 X46/X30/D0:neg DVDD:1031 0.866667
rDVDD/5569 X46/X30/D0:neg DVDD:1029 2.6
rDVDD/5570 X46/X30/D0:neg DVDD:954 5.2
rDVDD/5571 DVDD:945 DVDD:4190 0.0304865
rDVDD/5572 DVDD:945 X46/X30/D0:neg 1.73333
rDVDD/5573 DVDD:943 DVDD:4188 0.0571622
rDVDD/5574 DVDD:943 X46/X30/D0:neg 1.73333
rDVDD/5575 DVDD:941 DVDD:4186 0.0839189
rDVDD/5576 DVDD:941 DVDD:4183 2.25
rDVDD/5577 DVDD:941 DVDD:4168 0.0620347
rDVDD/5578 DVDD:941 X46/X30/D0:neg 0.866667
rDVDD/5579 DVDD:936 DVDD:4200 0.0304865
rDVDD/5580 DVDD:936 X46/X30/D0:neg 1.73333
rDVDD/5581 DVDD:934 DVDD:4198 0.0571622
rDVDD/5582 DVDD:934 X46/X30/D0:neg 1.73333
rDVDD/5583 DVDD:932 DVDD:4196 0.0839189
rDVDD/5584 DVDD:932 X46/X30/D0:neg 1.73333
rDVDD/5585 DVDD:929 DVDD:4210 0.0838378
rDVDD/5586 DVDD:929 X46/X30/D0:neg 1.73333
rDVDD/5587 DVDD:927 DVDD:4208 0.0570811
rDVDD/5588 DVDD:927 X46/X30/D0:neg 1.73333
rDVDD/5589 DVDD:925 DVDD:4206 0.0304054
rDVDD/5590 DVDD:925 X46/X30/D0:neg 1.73333
rDVDD/5591 DVDD:923 DVDD:4203 2.25
rDVDD/5592 DVDD:923 DVDD:4174 0.0945034
rDVDD/5593 DVDD:923 X46/X30/D0:neg 1.73333
rDVDD/5594 DVDD:920 DVDD:4220 0.0838378
rDVDD/5595 DVDD:920 X46/X30/D0:neg 1.73333
rDVDD/5596 DVDD:918 DVDD:4218 0.0570811
rDVDD/5597 DVDD:918 X46/X30/D0:neg 1.73333
rDVDD/5598 DVDD:916 DVDD:4216 0.0304054
rDVDD/5599 DVDD:916 X46/X30/D0:neg 1.73333
rDVDD/5600 DVDD:914 DVDD:4213 2.25
rDVDD/5601 DVDD:914 DVDD:4178 0.0945034
rDVDD/5602 DVDD:914 X46/X30/D0:neg 1.73333
rDVDD/5603 DVDD:911 DVDD:4004 0.00372973
rDVDD/5604 DVDD:911 X46/X30/D0:neg 1.73333
rDVDD/5605 DVDD:909 DVDD:4002 0.0304865
rDVDD/5606 DVDD:909 X46/X30/D0:neg 1.73333
rDVDD/5607 DVDD:907 DVDD:4000 0.0571622
rDVDD/5608 DVDD:907 X46/X30/D0:neg 1.73333
rDVDD/5609 DVDD:905 DVDD:3998 0.0839189
rDVDD/5610 DVDD:905 X46/X30/D0:neg 1.73333
rDVDD/5611 DVDD:902 DVDD:4014 0.00372973
rDVDD/5612 DVDD:902 X46/X30/D0:neg 1.73333
rDVDD/5613 DVDD:900 DVDD:4012 0.0304865
rDVDD/5614 DVDD:900 X46/X30/D0:neg 1.73333
rDVDD/5615 DVDD:898 DVDD:4010 0.0571622
rDVDD/5616 DVDD:898 X46/X30/D0:neg 1.73333
rDVDD/5617 DVDD:896 DVDD:4008 0.0839189
rDVDD/5618 DVDD:896 X46/X30/D0:neg 1.73333
rDVDD/5619 DVDD:893 DVDD:4024 0.00372973
rDVDD/5620 DVDD:893 DVDD:4022 0.0838378
rDVDD/5621 DVDD:893 X46/X30/D0:neg 1.73333
rDVDD/5622 DVDD:891 DVDD:4020 0.0570811
rDVDD/5623 DVDD:891 X46/X30/D0:neg 1.73333
rDVDD/5624 DVDD:889 DVDD:4018 0.0304054
rDVDD/5625 DVDD:889 X46/X30/D0:neg 1.73333
rDVDD/5626 DVDD:887 DVDD:4016 0.00364865
rDVDD/5627 DVDD:887 X46/X30/D0:neg 1.73333
rDVDD/5628 DVDD:884 DVDD:4034 0.00372973
rDVDD/5629 DVDD:884 DVDD:4032 0.0838378
rDVDD/5630 DVDD:884 X46/X30/D0:neg 1.73333
rDVDD/5631 DVDD:882 DVDD:4030 0.0570811
rDVDD/5632 DVDD:882 X46/X30/D0:neg 1.73333
rDVDD/5633 DVDD:880 DVDD:4028 0.0304054
rDVDD/5634 DVDD:880 X46/X30/D0:neg 1.73333
rDVDD/5635 DVDD:878 DVDD:4026 0.00364865
rDVDD/5636 DVDD:878 X46/X30/D0:neg 1.73333
rDVDD/5637 DVDD:875 DVDD:4222 8.10811e-05
rDVDD/5638 DVDD:875 DVDD:920 0.00364865
rDVDD/5639 DVDD:875 X46/X30/D0:neg 1.73333
rDVDD/5640 DVDD:873 DVDD:4220 0.0268378
rDVDD/5641 DVDD:873 DVDD:918 0.00364865
rDVDD/5642 DVDD:873 X46/X30/D0:neg 1.73333
rDVDD/5643 DVDD:871 DVDD:4218 0.0535946
rDVDD/5644 DVDD:871 DVDD:916 0.00356757
rDVDD/5645 DVDD:871 X46/X30/D0:neg 1.73333
rDVDD/5646 DVDD:869 DVDD:4216 0.0803514
rDVDD/5647 DVDD:869 DVDD:914 0.00356757
rDVDD/5648 DVDD:869 X46/X30/D0:neg 1.73333
rDVDD/5649 DVDD:865 DVDD:4212 0.00251351
rDVDD/5650 DVDD:865 DVDD:929 0.00121622
rDVDD/5651 DVDD:865 X46/X30/D0:neg 1.73333
rDVDD/5652 DVDD:863 DVDD:4210 0.0292703
rDVDD/5653 DVDD:863 DVDD:927 0.00121622
rDVDD/5654 DVDD:863 X46/X30/D0:neg 1.73333
rDVDD/5655 DVDD:861 DVDD:4208 0.056027
rDVDD/5656 DVDD:861 DVDD:925 0.00113514
rDVDD/5657 DVDD:861 X46/X30/D0:neg 1.73333
rDVDD/5658 DVDD:859 DVDD:4206 0.0827838
rDVDD/5659 DVDD:859 DVDD:923 0.00113514
rDVDD/5660 DVDD:859 X46/X30/D0:neg 1.73333
rDVDD/5661 DVDD:855 DVDD:4202 0.00486486
rDVDD/5662 DVDD:855 DVDD:4200 0.0827027
rDVDD/5663 DVDD:855 X46/X30/D0:neg 1.73333
rDVDD/5664 DVDD:853 DVDD:936 0.00113514
rDVDD/5665 DVDD:853 DVDD:4198 0.0559459
rDVDD/5666 DVDD:853 X46/X30/D0:neg 1.73333
rDVDD/5667 DVDD:851 DVDD:934 0.00121622
rDVDD/5668 DVDD:851 DVDD:4196 0.0291892
rDVDD/5669 DVDD:851 X46/X30/D0:neg 1.73333
rDVDD/5670 DVDD:849 DVDD:932 0.00121622
rDVDD/5671 DVDD:849 DVDD:4194 0.00243243
rDVDD/5672 DVDD:849 X46/X30/D0:neg 1.73333
rDVDD/5673 DVDD:845 DVDD:4192 0.0072973
rDVDD/5674 DVDD:845 DVDD:4190 0.0802703
rDVDD/5675 DVDD:845 X46/X30/D0:neg 1.73333
rDVDD/5676 DVDD:843 DVDD:945 0.00356757
rDVDD/5677 DVDD:843 DVDD:4188 0.0535135
rDVDD/5678 DVDD:843 X46/X30/D0:neg 1.73333
rDVDD/5679 DVDD:841 DVDD:943 0.00364865
rDVDD/5680 DVDD:841 DVDD:4186 0.0267568
rDVDD/5681 DVDD:841 X46/X30/D0:neg 1.73333
rDVDD/5682 DVDD:834 DVDD:4032 0.0268378
rDVDD/5683 DVDD:834 DVDD:882 0.00364865
rDVDD/5684 DVDD:834 X46/X30/D0:neg 1.73333
rDVDD/5685 DVDD:832 DVDD:4030 0.0535946
rDVDD/5686 DVDD:832 DVDD:880 0.00356757
rDVDD/5687 DVDD:832 X46/X30/D0:neg 1.73333
rDVDD/5688 DVDD:830 DVDD:4028 0.0803514
rDVDD/5689 DVDD:830 DVDD:878 0.00356757
rDVDD/5690 DVDD:830 X46/X30/D0:neg 1.73333
rDVDD/5691 DVDD:824 DVDD:4022 0.0292703
rDVDD/5692 DVDD:824 DVDD:891 0.00121622
rDVDD/5693 DVDD:824 X46/X30/D0:neg 1.73333
rDVDD/5694 DVDD:822 DVDD:4020 0.056027
rDVDD/5695 DVDD:822 DVDD:889 0.00113514
rDVDD/5696 DVDD:822 X46/X30/D0:neg 1.73333
rDVDD/5697 DVDD:820 DVDD:4018 0.0827838
rDVDD/5698 DVDD:820 DVDD:887 0.00113514
rDVDD/5699 DVDD:820 X46/X30/D0:neg 1.73333
rDVDD/5700 DVDD:816 DVDD:902 0.00113514
rDVDD/5701 DVDD:816 DVDD:4012 0.0827027
rDVDD/5702 DVDD:816 X46/X30/D0:neg 1.73333
rDVDD/5703 DVDD:814 DVDD:900 0.00113514
rDVDD/5704 DVDD:814 DVDD:4010 0.0559459
rDVDD/5705 DVDD:814 X46/X30/D0:neg 1.73333
rDVDD/5706 DVDD:812 DVDD:898 0.00121622
rDVDD/5707 DVDD:812 DVDD:4008 0.0291892
rDVDD/5708 DVDD:812 X46/X30/D0:neg 1.73333
rDVDD/5709 DVDD:810 DVDD:896 0.00121622
rDVDD/5710 DVDD:810 DVDD:4006 0.00243243
rDVDD/5711 DVDD:810 X46/X30/D0:neg 1.73333
rDVDD/5712 DVDD:806 DVDD:911 0.00356757
rDVDD/5713 DVDD:806 DVDD:4002 0.0802703
rDVDD/5714 DVDD:806 X46/X30/D0:neg 1.73333
rDVDD/5715 DVDD:804 DVDD:909 0.00356757
rDVDD/5716 DVDD:804 DVDD:4000 0.0535135
rDVDD/5717 DVDD:804 X46/X30/D0:neg 1.73333
rDVDD/5718 DVDD:802 DVDD:907 0.00364865
rDVDD/5719 DVDD:802 DVDD:3998 0.0267568
rDVDD/5720 DVDD:802 X46/X30/D0:neg 1.73333
rDVDD/5721 DVDD:800 DVDD:3995 2.25
rDVDD/5722 DVDD:800 DVDD:905 0.00364865
rDVDD/5723 DVDD:800 DVDD:3980 0.058386
rDVDD/5724 DVDD:800 X46/X30/D0:neg 1.73333
rDVDD/5725 DVDD:795 X46/D0:neg 0.67826
rDVDD/5726 DVDD:793 X46/D0:neg 0.67826
rDVDD/5727 DVDD:791 X46/D0:neg 0.67826
rDVDD/5728 DVDD:789 X46/D0:neg 0.67826
rDVDD/5729 DVDD:787 X46/D0:neg 0.67826
rDVDD/5730 DVDD:785 X46/D0:neg 0.67826
rDVDD/5731 DVDD:783 X46/D0:neg 0.67826
rDVDD/5732 DVDD:781 X46/D0:neg 0.67826
rDVDD/5733 DVDD:779 X46/D0:neg 0.67826
rDVDD/5734 DVDD:777 X46/D0:neg 0.67826
rDVDD/5735 DVDD:775 X46/D0:neg 0.67826
rDVDD/5736 DVDD:773 X46/D0:neg 0.67826
rDVDD/5737 DVDD:771 X46/D0:neg 0.67826
rDVDD/5738 DVDD:765 DVDD:795 0.0192308
rDVDD/5739 DVDD:765 X46/D0:neg 0.67826
rDVDD/5740 DVDD:763 DVDD:793 0.0192308
rDVDD/5741 DVDD:763 X46/D0:neg 0.67826
rDVDD/5742 DVDD:761 DVDD:791 0.0192308
rDVDD/5743 DVDD:761 X46/D0:neg 0.67826
rDVDD/5744 DVDD:759 DVDD:789 0.0192308
rDVDD/5745 DVDD:759 X46/D0:neg 0.67826
rDVDD/5746 DVDD:757 DVDD:787 0.0384615
rDVDD/5747 DVDD:757 X46/D0:neg 0.67826
rDVDD/5748 DVDD:755 DVDD:785 0.0192308
rDVDD/5749 DVDD:755 X46/D0:neg 0.67826
rDVDD/5750 DVDD:753 DVDD:783 0.0192308
rDVDD/5751 DVDD:753 X46/D0:neg 0.67826
rDVDD/5752 DVDD:751 DVDD:781 0.0192308
rDVDD/5753 DVDD:751 X46/D0:neg 0.67826
rDVDD/5754 DVDD:749 DVDD:779 0.0192308
rDVDD/5755 DVDD:749 X46/D0:neg 0.67826
rDVDD/5756 DVDD:747 DVDD:777 0.0384615
rDVDD/5757 DVDD:747 X46/D0:neg 0.67826
rDVDD/5758 DVDD:745 DVDD:775 0.0192308
rDVDD/5759 DVDD:745 X46/D0:neg 0.67826
rDVDD/5760 DVDD:743 DVDD:773 0.0192308
rDVDD/5761 DVDD:743 X46/D0:neg 0.67826
rDVDD/5762 DVDD:741 DVDD:771 0.0192308
rDVDD/5763 DVDD:741 X46/D0:neg 0.67826
rDVDD/5764 DVDD:735 DVDD:1943 0.0482197
rDVDD/5765 DVDD:735 DVDD:795 0.0378736
rDVDD/5766 DVDD:735 X46/D0:neg 0.226087
rDVDD/5767 DVDD:733 DVDD:765 0.0384615
rDVDD/5768 DVDD:733 DVDD:793 0.0384615
rDVDD/5769 DVDD:733 X46/D0:neg 0.67826
rDVDD/5770 DVDD:731 DVDD:763 0.0192308
rDVDD/5771 DVDD:731 DVDD:791 0.0384615
rDVDD/5772 DVDD:731 X46/D0:neg 0.67826
rDVDD/5773 DVDD:729 DVDD:761 0.0384615
rDVDD/5774 DVDD:729 DVDD:789 0.0384615
rDVDD/5775 DVDD:729 X46/D0:neg 0.67826
rDVDD/5776 DVDD:727 DVDD:759 0.0384615
rDVDD/5777 DVDD:727 DVDD:787 0.0192308
rDVDD/5778 DVDD:727 X46/D0:neg 0.67826
rDVDD/5779 DVDD:725 DVDD:757 0.0192308
rDVDD/5780 DVDD:725 DVDD:785 0.0384615
rDVDD/5781 DVDD:725 X46/D0:neg 0.67826
rDVDD/5782 DVDD:723 DVDD:755 0.0384615
rDVDD/5783 DVDD:723 DVDD:783 0.0384615
rDVDD/5784 DVDD:723 X46/D0:neg 0.67826
rDVDD/5785 DVDD:721 DVDD:753 0.0191923
rDVDD/5786 DVDD:721 DVDD:781 0.0384615
rDVDD/5787 DVDD:721 X46/D0:neg 0.67826
rDVDD/5788 DVDD:719 DVDD:751 0.0384615
rDVDD/5789 DVDD:719 DVDD:779 0.0384615
rDVDD/5790 DVDD:719 X46/D0:neg 0.67826
rDVDD/5791 DVDD:717 DVDD:749 0.0384615
rDVDD/5792 DVDD:717 DVDD:777 0.0192308
rDVDD/5793 DVDD:717 X46/D0:neg 0.67826
rDVDD/5794 DVDD:715 DVDD:747 0.0192308
rDVDD/5795 DVDD:715 DVDD:775 0.0384615
rDVDD/5796 DVDD:715 X46/D0:neg 0.67826
rDVDD/5797 DVDD:713 DVDD:745 0.0384615
rDVDD/5798 DVDD:713 DVDD:773 0.0384615
rDVDD/5799 DVDD:713 X46/D0:neg 0.67826
rDVDD/5800 DVDD:711 DVDD:743 0.0192308
rDVDD/5801 DVDD:711 DVDD:771 0.0384615
rDVDD/5802 DVDD:711 X46/D0:neg 0.67826
rDVDD/5803 DVDD:709 DVDD:741 0.0384615
rDVDD/5804 DVDD:709 X46/D0:neg 0.67826
rDVDD/5805 DVDD:707 DVDD:2096 0.0482197
rDVDD/5806 DVDD:707 DVDD:709 0.0570659
rDVDD/5807 DVDD:707 X46/D0:neg 0.185714
rDVDD/5808 DVDD:702 X46/D0:neg 0.67826
rDVDD/5809 DVDD:700 X46/D0:neg 0.67826
rDVDD/5810 DVDD:698 X46/D0:neg 0.67826
rDVDD/5811 DVDD:696 X46/D0:neg 0.67826
rDVDD/5812 DVDD:694 X46/D0:neg 0.67826
rDVDD/5813 DVDD:692 X46/D0:neg 0.67826
rDVDD/5814 DVDD:690 X46/D0:neg 0.67826
rDVDD/5815 DVDD:688 X46/D0:neg 0.67826
rDVDD/5816 DVDD:686 X46/D0:neg 0.67826
rDVDD/5817 DVDD:684 X46/D0:neg 0.67826
rDVDD/5818 DVDD:682 X46/D0:neg 0.67826
rDVDD/5819 DVDD:680 X46/D0:neg 0.67826
rDVDD/5820 DVDD:678 X46/D0:neg 0.67826
rDVDD/5821 DVDD:672 DVDD:702 0.0192308
rDVDD/5822 DVDD:672 X46/D0:neg 0.67826
rDVDD/5823 DVDD:670 DVDD:700 0.0192308
rDVDD/5824 DVDD:670 X46/D0:neg 0.67826
rDVDD/5825 DVDD:668 DVDD:698 0.0192308
rDVDD/5826 DVDD:668 X46/D0:neg 0.67826
rDVDD/5827 DVDD:666 DVDD:696 0.0192308
rDVDD/5828 DVDD:666 X46/D0:neg 0.67826
rDVDD/5829 DVDD:664 DVDD:694 0.0384615
rDVDD/5830 DVDD:664 X46/D0:neg 0.67826
rDVDD/5831 DVDD:662 DVDD:692 0.0192308
rDVDD/5832 DVDD:662 X46/D0:neg 0.67826
rDVDD/5833 DVDD:660 DVDD:690 0.0192308
rDVDD/5834 DVDD:660 X46/D0:neg 0.67826
rDVDD/5835 DVDD:658 DVDD:688 0.0192308
rDVDD/5836 DVDD:658 X46/D0:neg 0.67826
rDVDD/5837 DVDD:656 DVDD:686 0.0192308
rDVDD/5838 DVDD:656 X46/D0:neg 0.67826
rDVDD/5839 DVDD:654 DVDD:684 0.0384615
rDVDD/5840 DVDD:654 X46/D0:neg 0.67826
rDVDD/5841 DVDD:652 DVDD:682 0.0192308
rDVDD/5842 DVDD:652 X46/D0:neg 0.67826
rDVDD/5843 DVDD:650 DVDD:680 0.0192308
rDVDD/5844 DVDD:650 X46/D0:neg 0.67826
rDVDD/5845 DVDD:648 DVDD:678 0.0192308
rDVDD/5846 DVDD:648 X46/D0:neg 0.67826
rDVDD/5847 DVDD:642 DVDD:2093 0.0482582
rDVDD/5848 DVDD:642 DVDD:702 0.0378736
rDVDD/5849 DVDD:642 X46/D0:neg 0.226087
rDVDD/5850 DVDD:640 DVDD:672 0.0384615
rDVDD/5851 DVDD:640 DVDD:700 0.0384615
rDVDD/5852 DVDD:640 X46/D0:neg 0.67826
rDVDD/5853 DVDD:638 DVDD:670 0.0192308
rDVDD/5854 DVDD:638 DVDD:698 0.0384615
rDVDD/5855 DVDD:638 X46/D0:neg 0.67826
rDVDD/5856 DVDD:636 DVDD:668 0.0384615
rDVDD/5857 DVDD:636 DVDD:696 0.0384615
rDVDD/5858 DVDD:636 X46/D0:neg 0.67826
rDVDD/5859 DVDD:634 DVDD:666 0.0384615
rDVDD/5860 DVDD:634 DVDD:694 0.0192308
rDVDD/5861 DVDD:634 X46/D0:neg 0.67826
rDVDD/5862 DVDD:632 DVDD:664 0.0192308
rDVDD/5863 DVDD:632 DVDD:692 0.0384615
rDVDD/5864 DVDD:632 X46/D0:neg 0.67826
rDVDD/5865 DVDD:630 DVDD:662 0.0384615
rDVDD/5866 DVDD:630 DVDD:690 0.0384615
rDVDD/5867 DVDD:630 X46/D0:neg 0.67826
rDVDD/5868 DVDD:628 DVDD:660 0.0191923
rDVDD/5869 DVDD:628 DVDD:688 0.0384615
rDVDD/5870 DVDD:628 X46/D0:neg 0.67826
rDVDD/5871 DVDD:626 DVDD:658 0.0384615
rDVDD/5872 DVDD:626 DVDD:686 0.0384615
rDVDD/5873 DVDD:626 X46/D0:neg 0.67826
rDVDD/5874 DVDD:624 DVDD:656 0.0384615
rDVDD/5875 DVDD:624 DVDD:684 0.0192308
rDVDD/5876 DVDD:624 X46/D0:neg 0.67826
rDVDD/5877 DVDD:622 DVDD:654 0.0192308
rDVDD/5878 DVDD:622 DVDD:682 0.0384615
rDVDD/5879 DVDD:622 X46/D0:neg 0.67826
rDVDD/5880 DVDD:620 DVDD:652 0.0384615
rDVDD/5881 DVDD:620 DVDD:680 0.0384615
rDVDD/5882 DVDD:620 X46/D0:neg 0.67826
rDVDD/5883 DVDD:618 DVDD:650 0.0192308
rDVDD/5884 DVDD:618 DVDD:678 0.0384615
rDVDD/5885 DVDD:618 X46/D0:neg 0.67826
rDVDD/5886 DVDD:616 DVDD:648 0.0384615
rDVDD/5887 DVDD:616 X46/D0:neg 0.67826
rDVDD/5888 DVDD:614 DVDD:2246 0.0482582
rDVDD/5889 DVDD:614 DVDD:616 0.0570659
rDVDD/5890 DVDD:614 X46/D0:neg 0.185714
rDVDD/5891 DVDD:611 D8:neg 0.4
rDVDD/5892 DVDD:609 DVDD:611 0.0733696
rDVDD/5893 DVDD:609 D8:neg 0.4
rDVDD/5894 DVDD:607 DVDD:609 0.0733696
rDVDD/5895 DVDD:607 DVDD:12287 0.0322337
rDVDD/5896 DVDD:607 D8:neg 0.4
rDVDD/5897 DVDD:605 DVDD:12287 0.0411359
rDVDD/5898 DVDD:605 DVDD:12291 0.0116902
rDVDD/5899 DVDD:605 D8:neg 0.4
rDVDD/5900 DVDD:603 DVDD:12291 0.0861359
rDVDD/5901 DVDD:603 D8:neg 0.4
rDVDD/5902 DVDD:601 DVDD:603 0.0733696
rDVDD/5903 DVDD:601 D8:neg 0.4
rDVDD/5904 DVDD:599 DVDD:601 0.0733696
rDVDD/5905 DVDD:599 D8:neg 0.4
rDVDD/5906 DVDD:597 DVDD:599 0.0733696
rDVDD/5907 DVDD:597 D8:neg 0.4
rDVDD/5908 DVDD:595 DVDD:597 0.0978261
rDVDD/5909 DVDD:595 D8:neg 0.4
rDVDD/5910 DVDD:593 DVDD:595 0.0733696
rDVDD/5911 DVDD:593 DVDD:12300 0.0253859
rDVDD/5912 DVDD:593 D8:neg 0.4
rDVDD/5913 DVDD:591 DVDD:12300 0.0479837
rDVDD/5914 DVDD:591 DVDD:12304 0.00484239
rDVDD/5915 DVDD:591 D8:neg 0.4
rDVDD/5916 DVDD:589 DVDD:12304 0.0685272
rDVDD/5917 DVDD:589 D8:neg 0.4
rDVDD/5918 DVDD:587 DVDD:589 0.0978261
rDVDD/5919 DVDD:587 D8:neg 0.4
rDVDD/5920 DVDD:585 DVDD:587 0.0733696
rDVDD/5921 DVDD:585 D8:neg 0.4
rDVDD/5922 DVDD:583 DVDD:585 0.0733206
rDVDD/5923 DVDD:583 D8:neg 0.4
rDVDD/5924 DVDD:581 DVDD:583 0.0733696
rDVDD/5925 DVDD:581 D8:neg 0.4
rDVDD/5926 DVDD:579 DVDD:581 0.0978261
rDVDD/5927 DVDD:579 D8:neg 0.4
rDVDD/5928 DVDD:577 DVDD:579 0.0733696
rDVDD/5929 DVDD:577 DVDD:12314 0.0440217
rDVDD/5930 DVDD:577 D8:neg 0.4
rDVDD/5931 DVDD:575 DVDD:12314 0.0293478
rDVDD/5932 DVDD:575 DVDD:12318 0.0234783
rDVDD/5933 DVDD:575 D8:neg 0.4
rDVDD/5934 DVDD:573 DVDD:12318 0.0498913
rDVDD/5935 DVDD:573 D8:neg 0.4
rDVDD/5936 DVDD:571 DVDD:573 0.0978261
rDVDD/5937 DVDD:571 D8:neg 0.4
rDVDD/5938 DVDD:569 DVDD:571 0.0733696
rDVDD/5939 DVDD:569 D8:neg 0.4
rDVDD/5940 DVDD:567 DVDD:569 0.0733696
rDVDD/5941 DVDD:567 D8:neg 0.4
rDVDD/5942 DVDD:565 DVDD:567 0.0733696
rDVDD/5943 DVDD:565 D8:neg 0.4
rDVDD/5944 DVDD:563 DVDD:565 0.0978261
rDVDD/5945 DVDD:563 DVDD:12327 0.0371739
rDVDD/5946 DVDD:563 D8:neg 0.4
rDVDD/5947 DVDD:561 DVDD:12327 0.0361957
rDVDD/5948 DVDD:561 DVDD:12331 0.0166304
rDVDD/5949 DVDD:561 D8:neg 0.4
rDVDD/5950 DVDD:559 DVDD:12331 0.0567391
rDVDD/5951 DVDD:559 D8:neg 0.4
rDVDD/5952 DVDD:557 DVDD:559 0.0733696
rDVDD/5953 DVDD:557 D8:neg 0.4
rDVDD/5954 DVDD:555 DVDD:557 0.0733696
rDVDD/5955 DVDD:555 D8:neg 1.3
rDVDD/5956 DVDD:552 D8:neg 0.4
rDVDD/5957 DVDD:550 DVDD:552 0.0733696
rDVDD/5958 DVDD:550 D8:neg 0.4
rDVDD/5959 DVDD:548 DVDD:550 0.0733696
rDVDD/5960 DVDD:548 DVDD:12234 0.0322337
rDVDD/5961 DVDD:548 D8:neg 0.4
rDVDD/5962 DVDD:546 DVDD:12234 0.0411359
rDVDD/5963 DVDD:546 DVDD:12238 0.0116902
rDVDD/5964 DVDD:546 D8:neg 0.4
rDVDD/5965 DVDD:544 DVDD:12238 0.0861359
rDVDD/5966 DVDD:544 D8:neg 0.4
rDVDD/5967 DVDD:542 DVDD:544 0.0733696
rDVDD/5968 DVDD:542 D8:neg 0.4
rDVDD/5969 DVDD:540 DVDD:542 0.0733696
rDVDD/5970 DVDD:540 D8:neg 0.4
rDVDD/5971 DVDD:538 DVDD:540 0.0733696
rDVDD/5972 DVDD:538 D8:neg 0.4
rDVDD/5973 DVDD:536 DVDD:538 0.0978261
rDVDD/5974 DVDD:536 D8:neg 0.4
rDVDD/5975 DVDD:534 DVDD:536 0.0733696
rDVDD/5976 DVDD:534 DVDD:12247 0.0253859
rDVDD/5977 DVDD:534 D8:neg 0.4
rDVDD/5978 DVDD:532 DVDD:12247 0.0479837
rDVDD/5979 DVDD:532 DVDD:12251 0.00484239
rDVDD/5980 DVDD:532 D8:neg 0.4
rDVDD/5981 DVDD:530 DVDD:12251 0.0685272
rDVDD/5982 DVDD:530 D8:neg 0.4
rDVDD/5983 DVDD:528 DVDD:530 0.0978261
rDVDD/5984 DVDD:528 D8:neg 0.4
rDVDD/5985 DVDD:526 DVDD:528 0.0733696
rDVDD/5986 DVDD:526 D8:neg 0.4
rDVDD/5987 DVDD:524 DVDD:526 0.0733206
rDVDD/5988 DVDD:524 D8:neg 0.4
rDVDD/5989 DVDD:522 DVDD:524 0.0733696
rDVDD/5990 DVDD:522 D8:neg 0.4
rDVDD/5991 DVDD:520 DVDD:522 0.0978261
rDVDD/5992 DVDD:520 D8:neg 0.4
rDVDD/5993 DVDD:518 DVDD:520 0.0733696
rDVDD/5994 DVDD:518 DVDD:12261 0.0440217
rDVDD/5995 DVDD:518 D8:neg 0.4
rDVDD/5996 DVDD:516 DVDD:12261 0.0293478
rDVDD/5997 DVDD:516 DVDD:12265 0.0234783
rDVDD/5998 DVDD:516 D8:neg 0.4
rDVDD/5999 DVDD:514 DVDD:12265 0.0498913
rDVDD/6000 DVDD:514 D8:neg 0.4
rDVDD/6001 DVDD:512 DVDD:514 0.0978261
rDVDD/6002 DVDD:512 D8:neg 0.4
rDVDD/6003 DVDD:510 DVDD:512 0.0733696
rDVDD/6004 DVDD:510 D8:neg 0.4
rDVDD/6005 DVDD:508 DVDD:510 0.0733696
rDVDD/6006 DVDD:508 D8:neg 0.4
rDVDD/6007 DVDD:506 DVDD:508 0.0733696
rDVDD/6008 DVDD:506 D8:neg 0.4
rDVDD/6009 DVDD:504 DVDD:506 0.0978261
rDVDD/6010 DVDD:504 DVDD:12274 0.0371739
rDVDD/6011 DVDD:504 D8:neg 0.4
rDVDD/6012 DVDD:502 DVDD:12274 0.0361957
rDVDD/6013 DVDD:502 DVDD:12278 0.0166304
rDVDD/6014 DVDD:502 D8:neg 0.4
rDVDD/6015 DVDD:500 DVDD:12278 0.0567391
rDVDD/6016 DVDD:500 D8:neg 0.4
rDVDD/6017 DVDD:498 DVDD:500 0.0733696
rDVDD/6018 DVDD:498 D8:neg 0.4
rDVDD/6019 DVDD:496 DVDD:498 0.0733696
rDVDD/6020 DVDD:496 D8:neg 1.3
rDVDD/6021 X30/D0:neg DVDD:11884 1.73333
rDVDD/6022 X30/D0:neg DVDD:11881 1.73333
rDVDD/6023 X30/D0:neg DVDD:11878 1.73333
rDVDD/6024 X30/D0:neg DVDD:11875 1.73333
rDVDD/6025 X30/D0:neg DVDD:11852 1.73333
rDVDD/6026 X30/D0:neg DVDD:11849 1.73333
rDVDD/6027 X30/D0:neg DVDD:11823 0.894532
rDVDD/6028 X30/D0:neg DVDD:11910 1.31989
rDVDD/6029 DVDD:488 DVDD:11826 0.02565
rDVDD/6030 DVDD:488 X30/D0:neg 1.73333
rDVDD/6031 DVDD:486 DVDD:488 0.04545
rDVDD/6032 DVDD:486 DVDD:11831 0.0261
rDVDD/6033 DVDD:486 X30/D0:neg 1.73333
rDVDD/6034 DVDD:484 DVDD:11834 0.0162
rDVDD/6035 DVDD:484 X30/D0:neg 1.73333
rDVDD/6036 DVDD:482 DVDD:484 0.04545
rDVDD/6037 DVDD:482 X30/D0:neg 1.73333
rDVDD/6038 DVDD:480 DVDD:482 0.0909
rDVDD/6039 DVDD:480 X30/D0:neg 1.73333
rDVDD/6040 DVDD:478 DVDD:480 0.04545
rDVDD/6041 DVDD:478 X30/D0:neg 1.73333
rDVDD/6042 DVDD:476 DVDD:478 0.0909
rDVDD/6043 DVDD:476 X30/D0:neg 1.73333
rDVDD/6044 DVDD:474 DVDD:476 0.04545
rDVDD/6045 DVDD:474 X30/D0:neg 1.73333
rDVDD/6046 DVDD:472 DVDD:474 0.0909
rDVDD/6047 DVDD:472 X30/D0:neg 1.73333
rDVDD/6048 DVDD:470 DVDD:472 0.04545
rDVDD/6049 DVDD:470 X30/D0:neg 1.73333
rDVDD/6050 DVDD:468 DVDD:470 0.0909
rDVDD/6051 DVDD:468 X30/D0:neg 1.73333
rDVDD/6052 DVDD:466 DVDD:468 0.04545
rDVDD/6053 DVDD:466 X30/D0:neg 1.73333
rDVDD/6054 DVDD:464 DVDD:466 0.0909
rDVDD/6055 DVDD:464 X30/D0:neg 1.73333
rDVDD/6056 DVDD:462 DVDD:464 0.04545
rDVDD/6057 DVDD:462 DVDD:11849 0.0846
rDVDD/6058 DVDD:462 X30/D0:neg 1.73333
rDVDD/6059 DVDD:456 DVDD:11852 0.09405
rDVDD/6060 DVDD:456 DVDD:11850 1.5
rDVDD/6061 DVDD:456 X30/D0:neg 1.73333
rDVDD/6062 DVDD:454 DVDD:456 0.04545
rDVDD/6063 DVDD:454 DVDD:11853 4.5
rDVDD/6064 DVDD:454 X30/D0:neg 1.73333
rDVDD/6065 DVDD:452 DVDD:454 0.09
rDVDD/6066 DVDD:452 X30/D0:neg 1.73333
rDVDD/6067 DVDD:450 DVDD:452 0.045
rDVDD/6068 DVDD:450 X30/D0:neg 1.73333
rDVDD/6069 DVDD:448 DVDD:450 0.09
rDVDD/6070 DVDD:448 X30/D0:neg 1.73333
rDVDD/6071 DVDD:446 DVDD:448 0.045
rDVDD/6072 DVDD:446 X30/D0:neg 1.73333
rDVDD/6073 DVDD:444 DVDD:446 0.09
rDVDD/6074 DVDD:444 X30/D0:neg 1.73333
rDVDD/6075 DVDD:442 DVDD:444 0.045
rDVDD/6076 DVDD:442 X30/D0:neg 1.73333
rDVDD/6077 DVDD:440 DVDD:442 0.09
rDVDD/6078 DVDD:440 X30/D0:neg 1.73333
rDVDD/6079 DVDD:438 DVDD:440 0.045
rDVDD/6080 DVDD:438 X30/D0:neg 1.73333
rDVDD/6081 DVDD:436 DVDD:438 0.09
rDVDD/6082 DVDD:436 X30/D0:neg 1.73333
rDVDD/6083 DVDD:434 DVDD:436 0.045
rDVDD/6084 DVDD:434 X30/D0:neg 1.73333
rDVDD/6085 DVDD:432 DVDD:434 0.09
rDVDD/6086 DVDD:432 X30/D0:neg 1.73333
rDVDD/6087 DVDD:430 DVDD:432 0.045
rDVDD/6088 DVDD:430 X30/D0:neg 1.73333
rDVDD/6089 DVDD:428 DVDD:430 0.09
rDVDD/6090 DVDD:428 X30/D0:neg 1.73333
rDVDD/6091 DVDD:426 DVDD:428 0.045
rDVDD/6092 DVDD:426 DVDD:11875 0.0711
rDVDD/6093 DVDD:426 X30/D0:neg 1.73333
rDVDD/6094 DVDD:416 DVDD:11884 0.0945
rDVDD/6095 DVDD:416 X30/D0:neg 1.73333
rDVDD/6096 DVDD:414 DVDD:416 0.045
rDVDD/6097 DVDD:414 X30/D0:neg 1.73333
rDVDD/6098 DVDD:412 DVDD:414 0.09
rDVDD/6099 DVDD:412 X30/D0:neg 1.73333
rDVDD/6100 DVDD:410 DVDD:412 0.045
rDVDD/6101 DVDD:410 X30/D0:neg 1.73333
rDVDD/6102 DVDD:408 DVDD:410 0.09
rDVDD/6103 DVDD:408 X30/D0:neg 1.73333
rDVDD/6104 DVDD:406 DVDD:408 0.045
rDVDD/6105 DVDD:406 X30/D0:neg 1.73333
rDVDD/6106 DVDD:404 DVDD:406 0.09
rDVDD/6107 DVDD:404 X30/D0:neg 1.73333
rDVDD/6108 DVDD:402 DVDD:404 0.045
rDVDD/6109 DVDD:402 X30/D0:neg 1.73333
rDVDD/6110 DVDD:400 DVDD:402 0.09
rDVDD/6111 DVDD:400 X30/D0:neg 1.73333
rDVDD/6112 DVDD:398 DVDD:400 0.045
rDVDD/6113 DVDD:398 X30/D0:neg 1.73333
rDVDD/6114 DVDD:396 DVDD:398 0.09
rDVDD/6115 DVDD:396 X30/D0:neg 1.73333
rDVDD/6116 DVDD:394 DVDD:396 0.045
rDVDD/6117 DVDD:394 DVDD:11899 0.0135
rDVDD/6118 DVDD:394 X30/D0:neg 1.73333
rDVDD/6119 DVDD:392 DVDD:11902 0.0279
rDVDD/6120 DVDD:392 X30/D0:neg 1.73333
rDVDD/6121 DVDD:390 DVDD:392 0.045
rDVDD/6122 DVDD:390 DVDD:11907 0.0243
rDVDD/6123 DVDD:390 X30/D0:neg 1.73333
rDVDD/6124 X29/D0:neg DVDD:11788 1.73333
rDVDD/6125 X29/D0:neg DVDD:11785 1.73333
rDVDD/6126 X29/D0:neg DVDD:11782 1.73333
rDVDD/6127 X29/D0:neg DVDD:11779 1.73333
rDVDD/6128 X29/D0:neg DVDD:11756 1.73333
rDVDD/6129 X29/D0:neg DVDD:11753 1.73333
rDVDD/6130 X29/D0:neg DVDD:11727 0.894532
rDVDD/6131 X29/D0:neg DVDD:11814 1.31989
rDVDD/6132 DVDD:379 DVDD:11730 0.02565
rDVDD/6133 DVDD:379 X29/D0:neg 1.73333
rDVDD/6134 DVDD:377 DVDD:379 0.04545
rDVDD/6135 DVDD:377 DVDD:11735 0.0261
rDVDD/6136 DVDD:377 X29/D0:neg 1.73333
rDVDD/6137 DVDD:375 DVDD:11738 0.0162
rDVDD/6138 DVDD:375 X29/D0:neg 1.73333
rDVDD/6139 DVDD:373 DVDD:375 0.04545
rDVDD/6140 DVDD:373 X29/D0:neg 1.73333
rDVDD/6141 DVDD:371 DVDD:373 0.0909
rDVDD/6142 DVDD:371 X29/D0:neg 1.73333
rDVDD/6143 DVDD:369 DVDD:371 0.04545
rDVDD/6144 DVDD:369 X29/D0:neg 1.73333
rDVDD/6145 DVDD:367 DVDD:369 0.0909
rDVDD/6146 DVDD:367 X29/D0:neg 1.73333
rDVDD/6147 DVDD:365 DVDD:367 0.04545
rDVDD/6148 DVDD:365 X29/D0:neg 1.73333
rDVDD/6149 DVDD:363 DVDD:365 0.0909
rDVDD/6150 DVDD:363 X29/D0:neg 1.73333
rDVDD/6151 DVDD:361 DVDD:363 0.04545
rDVDD/6152 DVDD:361 X29/D0:neg 1.73333
rDVDD/6153 DVDD:359 DVDD:361 0.0909
rDVDD/6154 DVDD:359 X29/D0:neg 1.73333
rDVDD/6155 DVDD:357 DVDD:359 0.04545
rDVDD/6156 DVDD:357 X29/D0:neg 1.73333
rDVDD/6157 DVDD:355 DVDD:357 0.0909
rDVDD/6158 DVDD:355 X29/D0:neg 1.73333
rDVDD/6159 DVDD:353 DVDD:355 0.04545
rDVDD/6160 DVDD:353 DVDD:11753 0.0846
rDVDD/6161 DVDD:353 X29/D0:neg 1.73333
rDVDD/6162 DVDD:347 DVDD:11756 0.09405
rDVDD/6163 DVDD:347 DVDD:11754 1.5
rDVDD/6164 DVDD:347 X29/D0:neg 1.73333
rDVDD/6165 DVDD:345 DVDD:347 0.04545
rDVDD/6166 DVDD:345 DVDD:11757 4.5
rDVDD/6167 DVDD:345 X29/D0:neg 1.73333
rDVDD/6168 DVDD:343 DVDD:345 0.09
rDVDD/6169 DVDD:343 X29/D0:neg 1.73333
rDVDD/6170 DVDD:341 DVDD:343 0.045
rDVDD/6171 DVDD:341 X29/D0:neg 1.73333
rDVDD/6172 DVDD:339 DVDD:341 0.09
rDVDD/6173 DVDD:339 X29/D0:neg 1.73333
rDVDD/6174 DVDD:337 DVDD:339 0.045
rDVDD/6175 DVDD:337 X29/D0:neg 1.73333
rDVDD/6176 DVDD:335 DVDD:337 0.09
rDVDD/6177 DVDD:335 X29/D0:neg 1.73333
rDVDD/6178 DVDD:333 DVDD:335 0.045
rDVDD/6179 DVDD:333 X29/D0:neg 1.73333
rDVDD/6180 DVDD:331 DVDD:333 0.09
rDVDD/6181 DVDD:331 X29/D0:neg 1.73333
rDVDD/6182 DVDD:329 DVDD:331 0.045
rDVDD/6183 DVDD:329 X29/D0:neg 1.73333
rDVDD/6184 DVDD:327 DVDD:329 0.09
rDVDD/6185 DVDD:327 X29/D0:neg 1.73333
rDVDD/6186 DVDD:325 DVDD:327 0.045
rDVDD/6187 DVDD:325 X29/D0:neg 1.73333
rDVDD/6188 DVDD:323 DVDD:325 0.09
rDVDD/6189 DVDD:323 X29/D0:neg 1.73333
rDVDD/6190 DVDD:321 DVDD:323 0.045
rDVDD/6191 DVDD:321 X29/D0:neg 1.73333
rDVDD/6192 DVDD:319 DVDD:321 0.09
rDVDD/6193 DVDD:319 X29/D0:neg 1.73333
rDVDD/6194 DVDD:317 DVDD:319 0.045
rDVDD/6195 DVDD:317 DVDD:11779 0.0711
rDVDD/6196 DVDD:317 X29/D0:neg 1.73333
rDVDD/6197 DVDD:307 DVDD:11788 0.0945
rDVDD/6198 DVDD:307 X29/D0:neg 1.73333
rDVDD/6199 DVDD:305 DVDD:307 0.045
rDVDD/6200 DVDD:305 X29/D0:neg 1.73333
rDVDD/6201 DVDD:303 DVDD:305 0.09
rDVDD/6202 DVDD:303 X29/D0:neg 1.73333
rDVDD/6203 DVDD:301 DVDD:303 0.045
rDVDD/6204 DVDD:301 X29/D0:neg 1.73333
rDVDD/6205 DVDD:299 DVDD:301 0.09
rDVDD/6206 DVDD:299 X29/D0:neg 1.73333
rDVDD/6207 DVDD:297 DVDD:299 0.045
rDVDD/6208 DVDD:297 X29/D0:neg 1.73333
rDVDD/6209 DVDD:295 DVDD:297 0.09
rDVDD/6210 DVDD:295 X29/D0:neg 1.73333
rDVDD/6211 DVDD:293 DVDD:295 0.045
rDVDD/6212 DVDD:293 X29/D0:neg 1.73333
rDVDD/6213 DVDD:291 DVDD:293 0.09
rDVDD/6214 DVDD:291 X29/D0:neg 1.73333
rDVDD/6215 DVDD:289 DVDD:291 0.045
rDVDD/6216 DVDD:289 X29/D0:neg 1.73333
rDVDD/6217 DVDD:287 DVDD:289 0.09
rDVDD/6218 DVDD:287 X29/D0:neg 1.73333
rDVDD/6219 DVDD:285 DVDD:287 0.045
rDVDD/6220 DVDD:285 DVDD:11803 0.0135
rDVDD/6221 DVDD:285 X29/D0:neg 1.73333
rDVDD/6222 DVDD:283 DVDD:11806 0.0279
rDVDD/6223 DVDD:283 X29/D0:neg 1.73333
rDVDD/6224 DVDD:281 DVDD:283 0.045
rDVDD/6225 DVDD:281 DVDD:11811 0.0243
rDVDD/6226 DVDD:281 X29/D0:neg 1.73333
rDVDD/6227 X28/D0:neg DVDD:11692 1.73333
rDVDD/6228 X28/D0:neg DVDD:11689 1.73333
rDVDD/6229 X28/D0:neg DVDD:11686 1.73333
rDVDD/6230 X28/D0:neg DVDD:11683 1.73333
rDVDD/6231 X28/D0:neg DVDD:11660 1.73333
rDVDD/6232 X28/D0:neg DVDD:11657 1.73333
rDVDD/6233 X28/D0:neg DVDD:11631 0.894532
rDVDD/6234 X28/D0:neg DVDD:11718 1.31989
rDVDD/6235 DVDD:270 DVDD:11634 0.02565
rDVDD/6236 DVDD:270 X28/D0:neg 1.73333
rDVDD/6237 DVDD:268 DVDD:270 0.04545
rDVDD/6238 DVDD:268 DVDD:11639 0.0261
rDVDD/6239 DVDD:268 X28/D0:neg 1.73333
rDVDD/6240 DVDD:266 DVDD:11642 0.0162
rDVDD/6241 DVDD:266 X28/D0:neg 1.73333
rDVDD/6242 DVDD:264 DVDD:266 0.04545
rDVDD/6243 DVDD:264 X28/D0:neg 1.73333
rDVDD/6244 DVDD:262 DVDD:264 0.0909
rDVDD/6245 DVDD:262 X28/D0:neg 1.73333
rDVDD/6246 DVDD:260 DVDD:262 0.04545
rDVDD/6247 DVDD:260 X28/D0:neg 1.73333
rDVDD/6248 DVDD:258 DVDD:260 0.0909
rDVDD/6249 DVDD:258 X28/D0:neg 1.73333
rDVDD/6250 DVDD:256 DVDD:258 0.04545
rDVDD/6251 DVDD:256 X28/D0:neg 1.73333
rDVDD/6252 DVDD:254 DVDD:256 0.0909
rDVDD/6253 DVDD:254 X28/D0:neg 1.73333
rDVDD/6254 DVDD:252 DVDD:254 0.04545
rDVDD/6255 DVDD:252 X28/D0:neg 1.73333
rDVDD/6256 DVDD:250 DVDD:252 0.0909
rDVDD/6257 DVDD:250 X28/D0:neg 1.73333
rDVDD/6258 DVDD:248 DVDD:250 0.04545
rDVDD/6259 DVDD:248 X28/D0:neg 1.73333
rDVDD/6260 DVDD:246 DVDD:248 0.0909
rDVDD/6261 DVDD:246 X28/D0:neg 1.73333
rDVDD/6262 DVDD:244 DVDD:246 0.04545
rDVDD/6263 DVDD:244 DVDD:11657 0.0846
rDVDD/6264 DVDD:244 X28/D0:neg 1.73333
rDVDD/6265 DVDD:238 DVDD:11660 0.09405
rDVDD/6266 DVDD:238 DVDD:11658 1.5
rDVDD/6267 DVDD:238 X28/D0:neg 1.73333
rDVDD/6268 DVDD:236 DVDD:238 0.04545
rDVDD/6269 DVDD:236 DVDD:11661 4.5
rDVDD/6270 DVDD:236 X28/D0:neg 1.73333
rDVDD/6271 DVDD:234 DVDD:236 0.09
rDVDD/6272 DVDD:234 X28/D0:neg 1.73333
rDVDD/6273 DVDD:232 DVDD:234 0.045
rDVDD/6274 DVDD:232 X28/D0:neg 1.73333
rDVDD/6275 DVDD:230 DVDD:232 0.09
rDVDD/6276 DVDD:230 X28/D0:neg 1.73333
rDVDD/6277 DVDD:228 DVDD:230 0.045
rDVDD/6278 DVDD:228 X28/D0:neg 1.73333
rDVDD/6279 DVDD:226 DVDD:228 0.09
rDVDD/6280 DVDD:226 X28/D0:neg 1.73333
rDVDD/6281 DVDD:224 DVDD:226 0.045
rDVDD/6282 DVDD:224 X28/D0:neg 1.73333
rDVDD/6283 DVDD:222 DVDD:224 0.09
rDVDD/6284 DVDD:222 X28/D0:neg 1.73333
rDVDD/6285 DVDD:220 DVDD:222 0.045
rDVDD/6286 DVDD:220 X28/D0:neg 1.73333
rDVDD/6287 DVDD:218 DVDD:220 0.09
rDVDD/6288 DVDD:218 X28/D0:neg 1.73333
rDVDD/6289 DVDD:216 DVDD:218 0.045
rDVDD/6290 DVDD:216 X28/D0:neg 1.73333
rDVDD/6291 DVDD:214 DVDD:216 0.09
rDVDD/6292 DVDD:214 X28/D0:neg 1.73333
rDVDD/6293 DVDD:212 DVDD:214 0.045
rDVDD/6294 DVDD:212 X28/D0:neg 1.73333
rDVDD/6295 DVDD:210 DVDD:212 0.09
rDVDD/6296 DVDD:210 X28/D0:neg 1.73333
rDVDD/6297 DVDD:208 DVDD:210 0.045
rDVDD/6298 DVDD:208 DVDD:11683 0.0711
rDVDD/6299 DVDD:208 X28/D0:neg 1.73333
rDVDD/6300 DVDD:198 DVDD:11692 0.0945
rDVDD/6301 DVDD:198 X28/D0:neg 1.73333
rDVDD/6302 DVDD:196 DVDD:198 0.045
rDVDD/6303 DVDD:196 X28/D0:neg 1.73333
rDVDD/6304 DVDD:194 DVDD:196 0.09
rDVDD/6305 DVDD:194 X28/D0:neg 1.73333
rDVDD/6306 DVDD:192 DVDD:194 0.045
rDVDD/6307 DVDD:192 X28/D0:neg 1.73333
rDVDD/6308 DVDD:190 DVDD:192 0.09
rDVDD/6309 DVDD:190 X28/D0:neg 1.73333
rDVDD/6310 DVDD:188 DVDD:190 0.045
rDVDD/6311 DVDD:188 X28/D0:neg 1.73333
rDVDD/6312 DVDD:186 DVDD:188 0.09
rDVDD/6313 DVDD:186 X28/D0:neg 1.73333
rDVDD/6314 DVDD:184 DVDD:186 0.045
rDVDD/6315 DVDD:184 X28/D0:neg 1.73333
rDVDD/6316 DVDD:182 DVDD:184 0.09
rDVDD/6317 DVDD:182 X28/D0:neg 1.73333
rDVDD/6318 DVDD:180 DVDD:182 0.045
rDVDD/6319 DVDD:180 X28/D0:neg 1.73333
rDVDD/6320 DVDD:178 DVDD:180 0.09
rDVDD/6321 DVDD:178 X28/D0:neg 1.73333
rDVDD/6322 DVDD:176 DVDD:178 0.045
rDVDD/6323 DVDD:176 DVDD:11707 0.0135
rDVDD/6324 DVDD:176 X28/D0:neg 1.73333
rDVDD/6325 DVDD:174 DVDD:11710 0.0279
rDVDD/6326 DVDD:174 X28/D0:neg 1.73333
rDVDD/6327 DVDD:172 DVDD:174 0.045
rDVDD/6328 DVDD:172 DVDD:11715 0.0243
rDVDD/6329 DVDD:172 X28/D0:neg 1.73333
rDVDD/6330 X27/D0:neg DVDD:11596 1.73333
rDVDD/6331 X27/D0:neg DVDD:11593 1.73333
rDVDD/6332 X27/D0:neg DVDD:11590 1.73333
rDVDD/6333 X27/D0:neg DVDD:11587 1.73333
rDVDD/6334 X27/D0:neg DVDD:11564 1.73333
rDVDD/6335 X27/D0:neg DVDD:11561 1.73333
rDVDD/6336 X27/D0:neg DVDD:11535 0.894532
rDVDD/6337 X27/D0:neg DVDD:11622 1.31989
rDVDD/6338 DVDD:161 DVDD:11538 0.02565
rDVDD/6339 DVDD:161 X27/D0:neg 1.73333
rDVDD/6340 DVDD:159 DVDD:161 0.04545
rDVDD/6341 DVDD:159 DVDD:11543 0.0261
rDVDD/6342 DVDD:159 X27/D0:neg 1.73333
rDVDD/6343 DVDD:157 DVDD:11546 0.0162
rDVDD/6344 DVDD:157 X27/D0:neg 1.73333
rDVDD/6345 DVDD:155 DVDD:157 0.04545
rDVDD/6346 DVDD:155 X27/D0:neg 1.73333
rDVDD/6347 DVDD:153 DVDD:155 0.0909
rDVDD/6348 DVDD:153 X27/D0:neg 1.73333
rDVDD/6349 DVDD:151 DVDD:153 0.04545
rDVDD/6350 DVDD:151 X27/D0:neg 1.73333
rDVDD/6351 DVDD:149 DVDD:151 0.0909
rDVDD/6352 DVDD:149 X27/D0:neg 1.73333
rDVDD/6353 DVDD:147 DVDD:149 0.04545
rDVDD/6354 DVDD:147 X27/D0:neg 1.73333
rDVDD/6355 DVDD:145 DVDD:147 0.0909
rDVDD/6356 DVDD:145 X27/D0:neg 1.73333
rDVDD/6357 DVDD:143 DVDD:145 0.04545
rDVDD/6358 DVDD:143 X27/D0:neg 1.73333
rDVDD/6359 DVDD:141 DVDD:143 0.0909
rDVDD/6360 DVDD:141 X27/D0:neg 1.73333
rDVDD/6361 DVDD:139 DVDD:141 0.04545
rDVDD/6362 DVDD:139 X27/D0:neg 1.73333
rDVDD/6363 DVDD:137 DVDD:139 0.0909
rDVDD/6364 DVDD:137 X27/D0:neg 1.73333
rDVDD/6365 DVDD:135 DVDD:137 0.04545
rDVDD/6366 DVDD:135 DVDD:11561 0.0846
rDVDD/6367 DVDD:135 X27/D0:neg 1.73333
rDVDD/6368 DVDD:129 DVDD:11564 0.09405
rDVDD/6369 DVDD:129 DVDD:11562 1.5
rDVDD/6370 DVDD:129 X27/D0:neg 1.73333
rDVDD/6371 DVDD:127 DVDD:129 0.04545
rDVDD/6372 DVDD:127 DVDD:11565 4.5
rDVDD/6373 DVDD:127 X27/D0:neg 1.73333
rDVDD/6374 DVDD:125 DVDD:127 0.09
rDVDD/6375 DVDD:125 X27/D0:neg 1.73333
rDVDD/6376 DVDD:123 DVDD:125 0.045
rDVDD/6377 DVDD:123 X27/D0:neg 1.73333
rDVDD/6378 DVDD:121 DVDD:123 0.09
rDVDD/6379 DVDD:121 X27/D0:neg 1.73333
rDVDD/6380 DVDD:119 DVDD:121 0.045
rDVDD/6381 DVDD:119 X27/D0:neg 1.73333
rDVDD/6382 DVDD:117 DVDD:119 0.09
rDVDD/6383 DVDD:117 X27/D0:neg 1.73333
rDVDD/6384 DVDD:115 DVDD:117 0.045
rDVDD/6385 DVDD:115 X27/D0:neg 1.73333
rDVDD/6386 DVDD:113 DVDD:115 0.09
rDVDD/6387 DVDD:113 X27/D0:neg 1.73333
rDVDD/6388 DVDD:111 DVDD:113 0.045
rDVDD/6389 DVDD:111 X27/D0:neg 1.73333
rDVDD/6390 DVDD:109 DVDD:111 0.09
rDVDD/6391 DVDD:109 X27/D0:neg 1.73333
rDVDD/6392 DVDD:107 DVDD:109 0.045
rDVDD/6393 DVDD:107 X27/D0:neg 1.73333
rDVDD/6394 DVDD:105 DVDD:107 0.09
rDVDD/6395 DVDD:105 X27/D0:neg 1.73333
rDVDD/6396 DVDD:103 DVDD:105 0.045
rDVDD/6397 DVDD:103 X27/D0:neg 1.73333
rDVDD/6398 DVDD:101 DVDD:103 0.09
rDVDD/6399 DVDD:101 X27/D0:neg 1.73333
rDVDD/6400 DVDD:99 DVDD:101 0.045
rDVDD/6401 DVDD:99 DVDD:11587 0.0711
rDVDD/6402 DVDD:99 X27/D0:neg 1.73333
rDVDD/6403 DVDD:89 DVDD:11596 0.0945
rDVDD/6404 DVDD:89 X27/D0:neg 1.73333
rDVDD/6405 DVDD:87 DVDD:89 0.045
rDVDD/6406 DVDD:87 X27/D0:neg 1.73333
rDVDD/6407 DVDD:85 DVDD:87 0.09
rDVDD/6408 DVDD:85 X27/D0:neg 1.73333
rDVDD/6409 DVDD:83 DVDD:85 0.045
rDVDD/6410 DVDD:83 X27/D0:neg 1.73333
rDVDD/6411 DVDD:81 DVDD:83 0.09
rDVDD/6412 DVDD:81 X27/D0:neg 1.73333
rDVDD/6413 DVDD:79 DVDD:81 0.045
rDVDD/6414 DVDD:79 X27/D0:neg 1.73333
rDVDD/6415 DVDD:77 DVDD:79 0.09
rDVDD/6416 DVDD:77 X27/D0:neg 1.73333
rDVDD/6417 DVDD:75 DVDD:77 0.045
rDVDD/6418 DVDD:75 X27/D0:neg 1.73333
rDVDD/6419 DVDD:73 DVDD:75 0.09
rDVDD/6420 DVDD:73 X27/D0:neg 1.73333
rDVDD/6421 DVDD:71 DVDD:73 0.045
rDVDD/6422 DVDD:71 X27/D0:neg 1.73333
rDVDD/6423 DVDD:69 DVDD:71 0.09
rDVDD/6424 DVDD:69 X27/D0:neg 1.73333
rDVDD/6425 DVDD:67 DVDD:69 0.045
rDVDD/6426 DVDD:67 DVDD:11611 0.0135
rDVDD/6427 DVDD:67 X27/D0:neg 1.73333
rDVDD/6428 DVDD:65 DVDD:11614 0.0279
rDVDD/6429 DVDD:65 X27/D0:neg 1.73333
rDVDD/6430 DVDD:63 DVDD:65 0.045
rDVDD/6431 DVDD:63 DVDD:11619 0.0243
rDVDD/6432 DVDD:63 X27/D0:neg 1.73333
rDVDD/6433 DVDD:57 DVDD:496 0.0544906
rDVDD/6434 DVDD:57 D8:neg 0.371429
rDVDD/6435 DVDD:55 DVDD:57 0.041333
rDVDD/6436 DVDD:55 D8:neg 0.371429
rDVDD/6437 DVDD:53 DVDD:55 0.0978261
rDVDD/6438 DVDD:53 D8:neg 0.371429
rDVDD/6439 DVDD:51 DVDD:53 0.0733696
rDVDD/6440 DVDD:51 D8:neg 0.371429
rDVDD/6441 DVDD:49 DVDD:51 0.0978261
rDVDD/6442 DVDD:49 D8:neg 0.371429
rDVDD/6443 DVDD:47 DVDD:49 0.0733696
rDVDD/6444 DVDD:47 D8:neg 0.371429
rDVDD/6445 DVDD:45 DVDD:47 0.0978261
rDVDD/6446 DVDD:45 D8:neg 0.371429
rDVDD/6447 DVDD:43 DVDD:45 0.0733206
rDVDD/6448 DVDD:43 D8:neg 0.371429
rDVDD/6449 DVDD:41 DVDD:43 0.0978261
rDVDD/6450 DVDD:41 D8:neg 0.371429
rDVDD/6451 DVDD:39 DVDD:41 0.0733696
rDVDD/6452 DVDD:39 D8:neg 0.371429
rDVDD/6453 DVDD:37 DVDD:39 0.0978261
rDVDD/6454 DVDD:37 D8:neg 0.371429
rDVDD/6455 DVDD:35 DVDD:37 0.0733696
rDVDD/6456 DVDD:35 D8:neg 0.371429
rDVDD/6457 DVDD:33 DVDD:35 0.0978261
rDVDD/6458 DVDD:33 D8:neg 0.371429
rDVDD/6459 DVDD:31 DVDD:555 0.0544906
rDVDD/6460 DVDD:31 DVDD:33 0.0657406
rDVDD/6461 DVDD:31 D8:neg 0.371429
rDVDD/6462 DVDD:28 DVDD:552 0.0789961
rDVDD/6463 DVDD:28 D8:neg 0.371429
rDVDD/6464 DVDD:26 DVDD:28 0.041333
rDVDD/6465 DVDD:26 D8:neg 0.371429
rDVDD/6466 DVDD:24 DVDD:26 0.0978261
rDVDD/6467 DVDD:24 D8:neg 0.371429
rDVDD/6468 DVDD:22 DVDD:24 0.0733696
rDVDD/6469 DVDD:22 D8:neg 0.371429
rDVDD/6470 DVDD:20 DVDD:22 0.0978261
rDVDD/6471 DVDD:20 D8:neg 0.371429
rDVDD/6472 DVDD:18 DVDD:20 0.0733696
rDVDD/6473 DVDD:18 D8:neg 0.371429
rDVDD/6474 DVDD:16 DVDD:18 0.0978261
rDVDD/6475 DVDD:16 D8:neg 0.371429
rDVDD/6476 DVDD:14 DVDD:16 0.0733206
rDVDD/6477 DVDD:14 D8:neg 0.371429
rDVDD/6478 DVDD:12 DVDD:14 0.0978261
rDVDD/6479 DVDD:12 D8:neg 0.371429
rDVDD/6480 DVDD:10 DVDD:12 0.0733696
rDVDD/6481 DVDD:10 D8:neg 0.371429
rDVDD/6482 DVDD:8 DVDD:10 0.0978261
rDVDD/6483 DVDD:8 D8:neg 0.371429
rDVDD/6484 DVDD:6 DVDD:8 0.0733696
rDVDD/6485 DVDD:6 D8:neg 0.371429
rDVDD/6486 DVDD:4 DVDD:6 0.0978261
rDVDD/6487 DVDD:4 D8:neg 0.371429
rDVDD/6488 DVDD:2 DVDD:611 0.0789961
rDVDD/6489 DVDD:2 DVDD:4 0.0657406
rDVDD/6490 DVDD:2 D8:neg 0.371429
rDVDD/6491 X46/D1:neg X46/X30/D0:neg 0.01
rDVDD/6492 X46/X33/D0:neg X46/X30/D0:neg 0.01
rDVDD/6493 X46/X32/D0:neg X46/X30/D0:neg 0.01
rDVDD/6494 X46/X31/D0:neg X46/X30/D0:neg 0.01
cVDD/0 VDD:435 vss 66.3382f
cVDD/1 VDD:336 vss 28.0005f
cVDD/2 VDD:191 vss 19.5806f
cVDD/3 VDD:94 vss 19.5214f
rVDD/4 VDD:435 VDD:436 0.143617
rVDD/5 VDD:433 VDD:436 0.0365143
rVDD/6 VDD:432 VDD:435 0.0365143
rVDD/7 VDD:432 VDD:433 0.143617
rVDD/8 VDD:430 VDD:433 0.00912857
rVDD/9 VDD:429 VDD:432 0.00912857
rVDD/10 VDD:429 VDD:430 0.143617
rVDD/11 VDD:427 VDD:430 0.0456429
rVDD/12 VDD:426 VDD:429 0.0456429
rVDD/13 VDD:426 VDD:427 0.143617
rVDD/14 VDD:422 VDD:427 0.0365143
rVDD/15 VDD:421 VDD:426 0.0365143
rVDD/16 VDD:421 VDD:422 0.0718085
rVDD/17 VDD:419 VDD:422 0.0456429
rVDD/18 VDD:418 VDD:421 0.0456429
rVDD/19 VDD:418 VDD:419 0.143617
rVDD/20 VDD:413 VDD:418 0.0365143
rVDD/21 VDD:410 VDD:413 0.0456429
rVDD/22 VDD:405 VDD:410 0.0456429
rVDD/23 VDD:402 VDD:405 0.0456429
rVDD/24 VDD:397 VDD:402 0.0365143
rVDD/25 VDD:394 VDD:397 0.0456429
rVDD/26 VDD:391 VDD:394 0.0365143
rVDD/27 VDD:388 VDD:391 0.00912857
rVDD/28 VDD:385 VDD:388 0.0456429
rVDD/29 VDD:380 VDD:385 0.0365143
rVDD/30 VDD:380 VDD:381 0.0718085
rVDD/31 VDD:378 VDD:381 0.0456429
rVDD/32 VDD:377 VDD:380 0.0456429
rVDD/33 VDD:377 VDD:378 0.143617
rVDD/34 VDD:372 VDD:377 0.0365143
rVDD/35 VDD:369 VDD:372 0.0456429
rVDD/36 VDD:364 VDD:369 0.0456429
rVDD/37 VDD:361 VDD:364 0.0456429
rVDD/38 VDD:361 VDD:362 0.143617
rVDD/39 VDD:357 VDD 0.0438429
rVDD/40 VDD:357 VDD:362 0.0365143
rVDD/41 VDD:356 VDD:361 0.0365143
rVDD/42 VDD:356 VDD:357 0.0718085
rVDD/43 VDD:350 VDD 0.0018
rVDD/44 VDD:349 VDD 0.0018
rVDD/45 VDD:349 VDD:350 0.143617
rVDD/46 VDD:346 VDD:350 0.0365143
rVDD/47 VDD:346 VDD:349 0.180131
rVDD/48 VDD:336 VDD:337 0.143617
rVDD/49 VDD:334 VDD:337 0.0365143
rVDD/50 VDD:333 VDD:336 0.0365143
rVDD/51 VDD:333 VDD:334 0.143617
rVDD/52 VDD:331 VDD:334 0.00912857
rVDD/53 VDD:330 VDD:333 0.00912857
rVDD/54 VDD:330 VDD:331 0.143617
rVDD/55 VDD:328 VDD:331 0.0456429
rVDD/56 VDD:327 VDD:330 0.0456429
rVDD/57 VDD:327 VDD:328 0.143617
rVDD/58 VDD:323 VDD:328 0.0365143
rVDD/59 VDD:322 VDD:327 0.0365143
rVDD/60 VDD:322 VDD:323 0.0718085
rVDD/61 VDD:320 VDD:323 0.0456429
rVDD/62 VDD:319 VDD:322 0.0456429
rVDD/63 VDD:319 VDD:320 0.143617
rVDD/64 VDD:314 VDD:319 0.0365143
rVDD/65 VDD:311 VDD:314 0.0456429
rVDD/66 VDD:306 VDD:311 0.0456429
rVDD/67 VDD:303 VDD:306 0.0456429
rVDD/68 VDD:298 VDD:303 0.0365143
rVDD/69 VDD:295 VDD:298 0.0456429
rVDD/70 VDD:292 VDD:295 0.0365143
rVDD/71 VDD:289 VDD:292 0.00912857
rVDD/72 VDD:286 VDD:289 0.0456429
rVDD/73 VDD:281 VDD:286 0.0365143
rVDD/74 VDD:281 VDD:282 0.0718085
rVDD/75 VDD:279 VDD:282 0.0456429
rVDD/76 VDD:278 VDD:281 0.0456429
rVDD/77 VDD:278 VDD:279 0.143617
rVDD/78 VDD:273 VDD:278 0.0365143
rVDD/79 VDD:270 VDD:273 0.0456429
rVDD/80 VDD:265 VDD:270 0.0456429
rVDD/81 VDD:262 VDD:265 0.0456429
rVDD/82 VDD:262 VDD:263 0.143617
rVDD/83 VDD:258 VDD 0.0438429
rVDD/84 VDD:258 VDD:263 0.0365143
rVDD/85 VDD:257 VDD:262 0.0365143
rVDD/86 VDD:257 VDD:258 0.0718085
rVDD/87 VDD:251 VDD 0.0018
rVDD/88 VDD:250 VDD 0.0018
rVDD/89 VDD:250 VDD:251 0.143617
rVDD/90 VDD:247 VDD:251 0.0365143
rVDD/91 VDD:247 VDD:250 0.180131
rVDD/92 VDD:243 VDD:356 0.0327214
rVDD/93 VDD:239 VDD:243 4.5558
rVDD/94 VDD:236 VDD:239 0.0558
rVDD/95 VDD:233 VDD:236 0.1116
rVDD/96 VDD:230 VDD:233 0.0558
rVDD/97 VDD:227 VDD:230 0.1116
rVDD/98 VDD:224 VDD:227 0.0558
rVDD/99 VDD:222 VDD 0.00315
rVDD/100 VDD:222 VDD:239 1.5
rVDD/101 VDD:222 VDD:236 1.5
rVDD/102 VDD:222 VDD:233 1.5
rVDD/103 VDD:222 VDD:230 1.5
rVDD/104 VDD:222 VDD:227 1.5
rVDD/105 VDD:222 VDD:224 1.5
rVDD/106 VDD:222 VDD:243 0.00797143
rVDD/107 VDD:221 VDD:224 0.1116
rVDD/108 VDD:221 VDD:222 1.5
rVDD/109 VDD:219 VDD:257 0.0327214
rVDD/110 VDD:218 VDD:221 4.482
rVDD/111 VDD:218 VDD:219 4.5
rVDD/112 VDD:197 VDD 0.00315
rVDD/113 VDD:197 VDD:218 0.387402
rVDD/114 VDD:197 VDD:219 0.00797143
rVDD/115 VDD:191 VDD:435 0.166179
rVDD/116 VDD:191 VDD:436 0.0456429
rVDD/117 VDD:187 VDD:191 0.140821
rVDD/118 VDD:187 VDD:436 0.143617
rVDD/119 VDD:184 VDD:187 0.0162286
rVDD/120 VDD:184 VDD:433 0.143617
rVDD/121 VDD:181 VDD:184 0.00405714
rVDD/122 VDD:181 VDD:430 0.143617
rVDD/123 VDD:178 VDD:181 0.0202857
rVDD/124 VDD:178 VDD:427 0.143617
rVDD/125 VDD:173 VDD:178 0.0162286
rVDD/126 VDD:173 VDD:422 0.0718085
rVDD/127 VDD:170 VDD:173 0.0202857
rVDD/128 VDD:170 VDD:419 0.143617
rVDD/129 VDD:166 VDD:413 0.0718085
rVDD/130 VDD:166 VDD:419 0.0365143
rVDD/131 VDD:165 VDD:170 0.0162286
rVDD/132 VDD:165 VDD:166 0.0718085
rVDD/133 VDD:163 VDD:410 0.143617
rVDD/134 VDD:163 VDD:166 0.0456429
rVDD/135 VDD:162 VDD:165 0.0202857
rVDD/136 VDD:162 VDD:163 0.143617
rVDD/137 VDD:158 VDD:405 0.0718085
rVDD/138 VDD:158 VDD:163 0.0456429
rVDD/139 VDD:157 VDD:162 0.0202857
rVDD/140 VDD:157 VDD:158 0.0718085
rVDD/141 VDD:155 VDD:402 0.143617
rVDD/142 VDD:155 VDD:158 0.0456429
rVDD/143 VDD:154 VDD:157 0.0202857
rVDD/144 VDD:154 VDD:155 0.143617
rVDD/145 VDD:150 VDD:397 0.0718085
rVDD/146 VDD:150 VDD:155 0.0365143
rVDD/147 VDD:149 VDD:154 0.0162286
rVDD/148 VDD:149 VDD:150 0.0718085
rVDD/149 VDD:147 VDD:394 0.143617
rVDD/150 VDD:147 VDD:150 0.0456429
rVDD/151 VDD:146 VDD:149 0.0202857
rVDD/152 VDD:146 VDD:147 0.143617
rVDD/153 VDD:144 VDD:391 0.143617
rVDD/154 VDD:144 VDD:147 0.0365143
rVDD/155 VDD:143 VDD:146 0.0162286
rVDD/156 VDD:143 VDD:144 0.143617
rVDD/157 VDD:141 VDD:388 0.143617
rVDD/158 VDD:141 VDD:144 0.00912857
rVDD/159 VDD:140 VDD:143 0.00405714
rVDD/160 VDD:140 VDD:141 0.143617
rVDD/161 VDD:138 VDD:385 0.143617
rVDD/162 VDD:138 VDD:381 0.0365143
rVDD/163 VDD:138 VDD:141 0.0456429
rVDD/164 VDD:137 VDD:140 0.0202857
rVDD/165 VDD:137 VDD:138 0.143617
rVDD/166 VDD:132 VDD:137 0.0162286
rVDD/167 VDD:132 VDD:381 0.0718085
rVDD/168 VDD:129 VDD:132 0.0202857
rVDD/169 VDD:129 VDD:378 0.143617
rVDD/170 VDD:125 VDD:372 0.0718085
rVDD/171 VDD:125 VDD:378 0.0365143
rVDD/172 VDD:124 VDD:129 0.0162286
rVDD/173 VDD:124 VDD:125 0.0718085
rVDD/174 VDD:122 VDD:369 0.143617
rVDD/175 VDD:122 VDD:125 0.0456429
rVDD/176 VDD:121 VDD:124 0.0202857
rVDD/177 VDD:121 VDD:122 0.143617
rVDD/178 VDD:117 VDD:364 0.0718085
rVDD/179 VDD:117 VDD:362 0.0456429
rVDD/180 VDD:117 VDD:122 0.0456429
rVDD/181 VDD:116 VDD:121 0.0202857
rVDD/182 VDD:116 VDD:117 0.0718085
rVDD/183 VDD:113 VDD:116 0.0202857
rVDD/184 VDD:113 VDD:362 0.143617
rVDD/185 VDD:108 VDD:113 0.0162286
rVDD/186 VDD:108 VDD:357 0.0718085
rVDD/187 VDD VDD:108 0.0194857
rVDD/188 VDD:103 VDD 0.0008
rVDD/189 VDD:103 VDD:350 0.143617
rVDD/190 VDD:103 VDD:346 0.159846
rVDD/191 VDD:94 VDD:336 0.166179
rVDD/192 VDD:94 VDD:337 0.0456429
rVDD/193 VDD:90 VDD:94 0.140821
rVDD/194 VDD:90 VDD:337 0.143617
rVDD/195 VDD:87 VDD:90 0.0162286
rVDD/196 VDD:87 VDD:334 0.143617
rVDD/197 VDD:84 VDD:87 0.00405714
rVDD/198 VDD:84 VDD:331 0.143617
rVDD/199 VDD:81 VDD:84 0.0202857
rVDD/200 VDD:81 VDD:328 0.143617
rVDD/201 VDD:76 VDD:81 0.0162286
rVDD/202 VDD:76 VDD:323 0.0718085
rVDD/203 VDD:73 VDD:76 0.0202857
rVDD/204 VDD:73 VDD:320 0.143617
rVDD/205 VDD:69 VDD:314 0.0718085
rVDD/206 VDD:69 VDD:320 0.0365143
rVDD/207 VDD:68 VDD:73 0.0162286
rVDD/208 VDD:68 VDD:69 0.0718085
rVDD/209 VDD:66 VDD:311 0.143617
rVDD/210 VDD:66 VDD:69 0.0456429
rVDD/211 VDD:65 VDD:68 0.0202857
rVDD/212 VDD:65 VDD:66 0.143617
rVDD/213 VDD:61 VDD:306 0.0718085
rVDD/214 VDD:61 VDD:66 0.0456429
rVDD/215 VDD:60 VDD:65 0.0202857
rVDD/216 VDD:60 VDD:61 0.0718085
rVDD/217 VDD:58 VDD:303 0.143617
rVDD/218 VDD:58 VDD:61 0.0456429
rVDD/219 VDD:57 VDD:60 0.0202857
rVDD/220 VDD:57 VDD:58 0.143617
rVDD/221 VDD:53 VDD:298 0.0718085
rVDD/222 VDD:53 VDD:58 0.0365143
rVDD/223 VDD:52 VDD:57 0.0162286
rVDD/224 VDD:52 VDD:53 0.0718085
rVDD/225 VDD:50 VDD:295 0.143617
rVDD/226 VDD:50 VDD:53 0.0456429
rVDD/227 VDD:49 VDD:52 0.0202857
rVDD/228 VDD:49 VDD:50 0.143617
rVDD/229 VDD:47 VDD:292 0.143617
rVDD/230 VDD:47 VDD:50 0.0365143
rVDD/231 VDD:46 VDD:49 0.0162286
rVDD/232 VDD:46 VDD:47 0.143617
rVDD/233 VDD:44 VDD:289 0.143617
rVDD/234 VDD:44 VDD:47 0.00912857
rVDD/235 VDD:43 VDD:46 0.00405714
rVDD/236 VDD:43 VDD:44 0.143617
rVDD/237 VDD:41 VDD:286 0.143617
rVDD/238 VDD:41 VDD:282 0.0365143
rVDD/239 VDD:41 VDD:44 0.0456429
rVDD/240 VDD:40 VDD:43 0.0202857
rVDD/241 VDD:40 VDD:41 0.143617
rVDD/242 VDD:35 VDD:40 0.0162286
rVDD/243 VDD:35 VDD:282 0.0718085
rVDD/244 VDD:32 VDD:35 0.0202857
rVDD/245 VDD:32 VDD:279 0.143617
rVDD/246 VDD:28 VDD:273 0.0718085
rVDD/247 VDD:28 VDD:279 0.0365143
rVDD/248 VDD:27 VDD:32 0.0162286
rVDD/249 VDD:27 VDD:28 0.0718085
rVDD/250 VDD:25 VDD:270 0.143617
rVDD/251 VDD:25 VDD:28 0.0456429
rVDD/252 VDD:24 VDD:27 0.0202857
rVDD/253 VDD:24 VDD:25 0.143617
rVDD/254 VDD:20 VDD:265 0.0718085
rVDD/255 VDD:20 VDD:263 0.0456429
rVDD/256 VDD:20 VDD:25 0.0456429
rVDD/257 VDD:19 VDD:24 0.0202857
rVDD/258 VDD:19 VDD:20 0.0718085
rVDD/259 VDD:16 VDD:19 0.0202857
rVDD/260 VDD:16 VDD:263 0.143617
rVDD/261 VDD:11 VDD:16 0.0162286
rVDD/262 VDD:11 VDD:258 0.0718085
rVDD/263 VDD VDD:11 0.0194857
rVDD/264 VDD:6 VDD 0.0008
rVDD/265 VDD:6 VDD:251 0.143617
rVDD/266 VDD:6 VDD:247 0.159846
cPAD/0 PAD:15142 vss 0.500352f
cPAD/1 PAD:15004 vss 0.655995f
cPAD/2 PAD:14602 vss 0.533546f
cPAD/3 PAD:14601 vss 1.76086f
cPAD/4 PAD:9454 vss 0.533557f
cPAD/5 PAD:9453 vss 1.76087f
cPAD/6 PAD:9449 vss 0.23336f
cPAD/7 PAD:9304 vss 0.947604f
cPAD/8 PAD:8893 vss 13.2863f
cPAD/9 PAD:8891 vss 8.24412f
cPAD/10 PAD:8890 vss 3.62466f
cPAD/11 PAD:8723 vss 1.97215f
cPAD/12 PAD:8553 vss 1.52711f
cPAD/13 PAD:8383 vss 1.52711f
cPAD/14 PAD:8213 vss 1.52711f
cPAD/15 PAD:8043 vss 1.52711f
cPAD/16 PAD:7873 vss 1.52711f
cPAD/17 PAD:7703 vss 1.52711f
cPAD/18 PAD:7533 vss 1.52711f
cPAD/19 PAD:7363 vss 1.52711f
cPAD/20 PAD:7193 vss 1.52711f
cPAD/21 PAD:7023 vss 1.52711f
cPAD/22 PAD:6853 vss 1.52711f
cPAD/23 PAD:6683 vss 1.52711f
cPAD/24 PAD:6513 vss 1.52711f
cPAD/25 PAD:6343 vss 1.52711f
cPAD/26 PAD:6173 vss 1.52711f
cPAD/27 PAD:6003 vss 1.52711f
cPAD/28 PAD:5833 vss 1.52711f
cPAD/29 PAD:5663 vss 1.52711f
cPAD/30 PAD:5493 vss 1.52711f
cPAD/31 PAD:5323 vss 1.52711f
cPAD/32 PAD:5153 vss 1.52711f
cPAD/33 PAD:4983 vss 1.52711f
cPAD/34 PAD:4813 vss 1.52711f
cPAD/35 PAD:4643 vss 1.52711f
cPAD/36 PAD:4473 vss 1.52711f
cPAD/37 PAD:4303 vss 1.52711f
cPAD/38 PAD:4133 vss 1.52711f
cPAD/39 PAD:3963 vss 2.00416f
cPAD/40 PAD:3769 vss 5.61282f
cPAD/41 PAD:3725 vss 5.31154f
cPAD/42 R7:pos vss 0.072827f
cPAD/43 R6:pos vss 0.072827f
cPAD/44 R5:pos vss 0.072827f
cPAD/45 R4:pos vss 0.072827f
cPAD/46 R3:pos vss 0.072827f
rPAD/47 PAD:16978 PAD:16979 0.0786026
rPAD/48 PAD:15142 PAD:16890 0.0292349
rPAD/49 PAD:15137 PAD:16890 0.000724832
rPAD/50 PAD:15134 PAD:16832 0.0314094
rPAD/51 PAD:15134 PAD:15137 0.0599195
rPAD/52 PAD:15130 PAD:16774 0.0347919
rPAD/53 PAD:15130 PAD:16832 0.0135302
rPAD/54 PAD:15129 PAD:15130 0.346154
rPAD/55 PAD:15126 PAD:16716 0.0381745
rPAD/56 PAD:15126 PAD:16774 0.0101477
rPAD/57 PAD:15125 PAD:15126 0.346154
rPAD/58 PAD:15090 PAD:16194 0.0386577
rPAD/59 PAD:15090 PAD:16252 0.00966443
rPAD/60 PAD:15086 PAD:16136 0.0270604
rPAD/61 PAD:15086 PAD:16194 0.0212617
rPAD/62 PAD:15082 PAD:16078 0.030443
rPAD/63 PAD:15082 PAD:16136 0.0178792
rPAD/64 PAD:15038 PAD:15440 0.0227114
rPAD/65 PAD:15038 PAD:15498 0.0256107
rPAD/66 PAD:15034 PAD:15382 0.026094
rPAD/67 PAD:15034 PAD:15440 0.0222282
rPAD/68 PAD:15030 PAD:15324 0.0294765
rPAD/69 PAD:15030 PAD:15382 0.0188456
rPAD/70 PAD:15026 PAD:15266 0.0328591
rPAD/71 PAD:15026 PAD:15324 0.0154631
rPAD/72 PAD:15014 PAD:15017 0.0449396
rPAD/73 PAD:14987 PAD:14989 0.0182751
rPAD/74 PAD:14981 PAD:14983 0.0233843
rPAD/75 PAD:14971 PAD:14973 0.00569869
rPAD/76 PAD:14968 PAD:14971 0.0558079
rPAD/77 PAD:14966 PAD:14968 0.0170961
rPAD/78 PAD:14961 PAD:14963 0.0119869
rPAD/79 PAD:14948 PAD:17001 0.0524672
rPAD/80 PAD:14948 PAD:17003 0.0261354
rPAD/81 PAD:14947 PAD:14949 0.0261354
rPAD/82 PAD:14947 PAD:14948 0.9
rPAD/83 PAD:14945 PAD:14947 0.0524672
rPAD/84 PAD:14943 PAD:16999 0.0473581
rPAD/85 PAD:14943 PAD:17001 0.0312445
rPAD/86 PAD:14942 PAD:14943 0.9
rPAD/87 PAD:14940 PAD:14942 0.0473581
rPAD/88 PAD:14939 PAD:16997 0.0701528
rPAD/89 PAD:14939 PAD:16999 0.00844978
rPAD/90 PAD:14938 PAD:14940 0.00844978
rPAD/91 PAD:14938 PAD:14939 0.9
rPAD/92 PAD:14934 PAD:16997 0.013559
rPAD/93 PAD:14933 PAD:14935 0.013559
rPAD/94 PAD:14933 PAD:14934 0.9
rPAD/95 PAD:14930 PAD:16994 0.00923581
rPAD/96 PAD:14930 PAD:14934 0.0558079
rPAD/97 PAD:14929 PAD:14930 0.9
rPAD/98 PAD:14927 PAD:14929 0.00923581
rPAD/99 PAD:14924 PAD:16992 0.00412664
rPAD/100 PAD:14924 PAD:16994 0.074476
rPAD/101 PAD:14923 PAD:14924 0.9
rPAD/102 PAD:14921 PAD:14923 0.00412664
rPAD/103 PAD:14911 PAD:14913 0.0218122
rPAD/104 PAD:14909 PAD:14911 0.0339956
rPAD/105 PAD:14904 PAD:14906 0.0391048
rPAD/106 PAD:14899 PAD:14901 0.01631
rPAD/107 PAD:14893 PAD:14895 0.0214192
rPAD/108 PAD:14890 PAD:16979 0.00137555
rPAD/109 PAD:14889 PAD:14890 0.9
rPAD/110 PAD:14887 PAD:14889 0.00137555
rPAD/111 PAD:14884 PAD:16978 0.00373362
rPAD/112 PAD:14883 PAD:14885 0.00373362
rPAD/113 PAD:14883 PAD:14884 0.9
rPAD/114 PAD:14880 PAD:14883 0.0558079
rPAD/115 PAD:14878 PAD:14880 0.0190611
rPAD/116 PAD:14873 PAD:14875 0.013952
rPAD/117 PAD:14865 PAD:16969 0.0316376
rPAD/118 PAD:14865 PAD:16971 0.0469651
rPAD/119 PAD:14864 PAD:14865 0.9
rPAD/120 PAD:14860 PAD:16967 0.0544323
rPAD/121 PAD:14860 PAD:16969 0.0241703
rPAD/122 PAD:14855 PAD:16965 0.0493231
rPAD/123 PAD:14855 PAD:16967 0.0292795
rPAD/124 PAD:14850 PAD:14852 0.00648472
rPAD/125 PAD:14846 PAD:16963 0.0115939
rPAD/126 PAD:14845 PAD:14847 0.0115939
rPAD/127 PAD:14845 PAD:14846 0.9
rPAD/128 PAD:14842 PAD:16960 0.0112009
rPAD/129 PAD:14842 PAD:14846 0.0558079
rPAD/130 PAD:14841 PAD:14842 0.9
rPAD/131 PAD:14839 PAD:14841 0.0112009
rPAD/132 PAD:14836 PAD:16958 0.0060917
rPAD/133 PAD:14836 PAD:16960 0.0725109
rPAD/134 PAD:14835 PAD:14836 0.9
rPAD/135 PAD:14833 PAD:14835 0.0060917
rPAD/136 PAD:14831 PAD:16958 0.0497162
rPAD/137 PAD:14827 PAD:15144 0.0224017
rPAD/138 PAD:14827 PAD:14831 0.0925546
rPAD/139 PAD:14823 PAD:15144 0.00196507
rPAD/140 PAD:14822 PAD:14823 0.9
rPAD/141 PAD:14814 PAD:16890 0.026775
rPAD/142 PAD:14811 PAD:14814 0.0279
rPAD/143 PAD:14803 PAD:14806 0.01395
rPAD/144 PAD:14792 PAD:14795 0.01395
rPAD/145 PAD:14792 PAD:14793 0.586956
rPAD/146 PAD:14785 PAD:14788 0.01395
rPAD/147 PAD:14785 PAD:14786 0.586956
rPAD/148 PAD:14782 PAD:14785 0.01395
rPAD/149 PAD:14778 PAD:14779 0.586956
rPAD/150 PAD:14771 PAD:14774 0.01395
rPAD/151 PAD:14764 PAD:14767 0.01395
rPAD/152 PAD:14764 PAD:14765 0.586956
rPAD/153 PAD:14761 PAD:14765 0.0279
rPAD/154 PAD:14760 PAD:14761 0.586956
rPAD/155 PAD:14758 PAD:14761 0.01395
rPAD/156 PAD:14754 PAD:14758 0.0279
rPAD/157 PAD:14753 PAD:14754 0.586956
rPAD/158 PAD:14751 PAD:14754 0.01395
rPAD/159 PAD:14750 PAD:14753 0.01395
rPAD/160 PAD:14750 PAD:14751 0.586956
rPAD/161 PAD:14747 PAD:14751 0.0279
rPAD/162 PAD:14746 PAD:14747 0.586956
rPAD/163 PAD:14739 PAD:14742 0.01395
rPAD/164 PAD:14735 PAD:14736 0.586956
rPAD/165 PAD:14732 PAD:14735 0.01395
rPAD/166 PAD:14729 PAD:14732 0.01395
rPAD/167 PAD:14721 PAD:14722 0.586956
rPAD/168 PAD:14718 PAD:14721 0.01395
rPAD/169 PAD:14711 PAD:14714 0.01395
rPAD/170 PAD:14711 PAD:14712 0.586956
rPAD/171 PAD:14697 PAD:14700 0.01395
rPAD/172 PAD:14693 PAD:14694 0.586956
rPAD/173 PAD:14690 PAD:14694 0.0279
rPAD/174 PAD:14689 PAD:14690 0.586956
rPAD/175 PAD:14686 PAD:14689 0.01395
rPAD/176 PAD:14682 PAD:14683 0.586956
rPAD/177 PAD:14679 PAD:14682 0.01395
rPAD/178 PAD:14676 PAD:14679 0.01395
rPAD/179 PAD:14672 PAD:14673 0.586956
rPAD/180 PAD:14665 PAD:14668 0.01395
rPAD/181 PAD:14658 PAD:14661 0.01395
rPAD/182 PAD:14658 PAD:14659 0.586956
rPAD/183 PAD:14647 PAD:14648 0.586956
rPAD/184 PAD:14644 PAD:14647 0.01395
rPAD/185 PAD:14633 PAD:14636 0.01395
rPAD/186 PAD:14633 PAD:14634 0.586956
rPAD/187 PAD:14626 PAD:14629 0.01395
rPAD/188 PAD:14623 PAD:14626 0.01395
rPAD/189 PAD:14623 PAD:14624 0.586956
rPAD/190 PAD:14620 PAD:14624 0.0279
rPAD/191 PAD:14619 PAD:14620 0.586956
rPAD/192 PAD:14612 PAD:14615 0.01395
rPAD/193 PAD:14612 PAD:14613 0.586956
rPAD/194 PAD:14605 PAD:14608 0.01395
rPAD/195 PAD:14605 PAD:14606 0.586956
rPAD/196 PAD:14602 PAD:16889 0.01035
rPAD/197 PAD:14602 PAD:14606 0.0279
rPAD/198 PAD:14601 PAD:14602 0.586956
rPAD/199 PAD:14598 PAD:15000 0.000393013
rPAD/200 PAD:14598 PAD:14601 0.01035
rPAD/201 PAD:14597 PAD:16832 0.0100588
rPAD/202 PAD:14594 PAD:14597 0.0751765
rPAD/203 PAD:14591 PAD:14594 0.0375882
rPAD/204 PAD:14582 PAD:14585 0.0751765
rPAD/205 PAD:14579 PAD:14582 0.0375882
rPAD/206 PAD:14576 PAD:14579 0.0751765
rPAD/207 PAD:14573 PAD:14576 0.0375882
rPAD/208 PAD:14570 PAD:14573 0.0751765
rPAD/209 PAD:14567 PAD:14570 0.0375882
rPAD/210 PAD:14564 PAD:14567 0.0751765
rPAD/211 PAD:14561 PAD:14564 0.0375882
rPAD/212 PAD:14558 PAD:14561 0.0751765
rPAD/213 PAD:14555 PAD:14558 0.0375882
rPAD/214 PAD:14542 PAD:14545 0.0375882
rPAD/215 PAD:14539 PAD:14542 0.0751765
rPAD/216 PAD:14530 PAD:14533 0.0375882
rPAD/217 PAD:14525 PAD:14528 0.0375882
rPAD/218 PAD:14522 PAD:14525 0.0751765
rPAD/219 PAD:14519 PAD:14522 0.0375882
rPAD/220 PAD:14516 PAD:14519 0.0751765
rPAD/221 PAD:14513 PAD:14516 0.0375882
rPAD/222 PAD:14504 PAD:14507 0.0751765
rPAD/223 PAD:14501 PAD:14504 0.0375882
rPAD/224 PAD:14494 PAD:14497 0.0375882
rPAD/225 PAD:14491 PAD:14494 0.0751765
rPAD/226 PAD:14488 PAD:14491 0.0375882
rPAD/227 PAD:14485 PAD:14488 0.0751765
rPAD/228 PAD:14480 PAD:14483 0.0751765
rPAD/229 PAD:14471 PAD:14474 0.0375882
rPAD/230 PAD:14468 PAD:14471 0.0751765
rPAD/231 PAD:14465 PAD:14468 0.0375882
rPAD/232 PAD:14462 PAD:14465 0.0751765
rPAD/233 PAD:14459 PAD:14462 0.0375882
rPAD/234 PAD:14450 PAD:14453 0.0751765
rPAD/235 PAD:14447 PAD:14450 0.0375882
rPAD/236 PAD:14444 PAD:14447 0.0751765
rPAD/237 PAD:14441 PAD:14444 0.0375882
rPAD/238 PAD:14438 PAD:14441 0.0751765
rPAD/239 PAD:14435 PAD:14438 0.0375882
rPAD/240 PAD:14432 PAD:17018 0.0283817
rPAD/241 PAD:14432 PAD:14435 0.0751765
rPAD/242 PAD:14429 PAD:15129 0.0135302
rPAD/243 PAD:14427 PAD:16774 0.0100588
rPAD/244 PAD:14424 PAD:14427 0.0751765
rPAD/245 PAD:14421 PAD:14424 0.0375882
rPAD/246 PAD:14412 PAD:14415 0.0751765
rPAD/247 PAD:14409 PAD:14412 0.0375882
rPAD/248 PAD:14406 PAD:14409 0.0751765
rPAD/249 PAD:14403 PAD:14406 0.0375882
rPAD/250 PAD:14400 PAD:14403 0.0751765
rPAD/251 PAD:14397 PAD:14400 0.0375882
rPAD/252 PAD:14394 PAD:14397 0.0751765
rPAD/253 PAD:14391 PAD:14394 0.0375882
rPAD/254 PAD:14388 PAD:14391 0.0751765
rPAD/255 PAD:14385 PAD:14388 0.0375882
rPAD/256 PAD:14372 PAD:14375 0.0375882
rPAD/257 PAD:14369 PAD:14372 0.0751765
rPAD/258 PAD:14360 PAD:14363 0.0375882
rPAD/259 PAD:14355 PAD:14358 0.0375882
rPAD/260 PAD:14352 PAD:14355 0.0751765
rPAD/261 PAD:14349 PAD:14352 0.0375882
rPAD/262 PAD:14346 PAD:14349 0.0751765
rPAD/263 PAD:14343 PAD:14346 0.0375882
rPAD/264 PAD:14334 PAD:14337 0.0751765
rPAD/265 PAD:14331 PAD:14334 0.0375882
rPAD/266 PAD:14324 PAD:14327 0.0375882
rPAD/267 PAD:14321 PAD:14324 0.0751765
rPAD/268 PAD:14318 PAD:14321 0.0375882
rPAD/269 PAD:14315 PAD:14318 0.0751765
rPAD/270 PAD:14310 PAD:14313 0.0751765
rPAD/271 PAD:14301 PAD:14304 0.0375882
rPAD/272 PAD:14298 PAD:14301 0.0751765
rPAD/273 PAD:14295 PAD:14298 0.0375882
rPAD/274 PAD:14292 PAD:14295 0.0751765
rPAD/275 PAD:14289 PAD:14292 0.0375882
rPAD/276 PAD:14280 PAD:14283 0.0751765
rPAD/277 PAD:14277 PAD:14280 0.0375882
rPAD/278 PAD:14274 PAD:14277 0.0751765
rPAD/279 PAD:14271 PAD:14274 0.0375882
rPAD/280 PAD:14268 PAD:14271 0.0751765
rPAD/281 PAD:14265 PAD:14268 0.0375882
rPAD/282 PAD:14262 PAD:17016 0.0283817
rPAD/283 PAD:14262 PAD:14265 0.0751765
rPAD/284 PAD:14259 PAD:15125 0.0101477
rPAD/285 PAD:14259 PAD:15129 0.0347919
rPAD/286 PAD:14257 PAD:16716 0.0100588
rPAD/287 PAD:14254 PAD:14257 0.0751765
rPAD/288 PAD:14251 PAD:14254 0.0375882
rPAD/289 PAD:14242 PAD:14245 0.0751765
rPAD/290 PAD:14239 PAD:14242 0.0375882
rPAD/291 PAD:14236 PAD:14239 0.0751765
rPAD/292 PAD:14233 PAD:14236 0.0375882
rPAD/293 PAD:14230 PAD:14233 0.0751765
rPAD/294 PAD:14227 PAD:14230 0.0375882
rPAD/295 PAD:14224 PAD:14227 0.0751765
rPAD/296 PAD:14221 PAD:14224 0.0375882
rPAD/297 PAD:14218 PAD:14221 0.0751765
rPAD/298 PAD:14215 PAD:14218 0.0375882
rPAD/299 PAD:14202 PAD:14205 0.0375882
rPAD/300 PAD:14199 PAD:14202 0.0751765
rPAD/301 PAD:14190 PAD:14193 0.0375882
rPAD/302 PAD:14185 PAD:14188 0.0375882
rPAD/303 PAD:14182 PAD:14185 0.0751765
rPAD/304 PAD:14179 PAD:14182 0.0375882
rPAD/305 PAD:14176 PAD:14179 0.0751765
rPAD/306 PAD:14173 PAD:14176 0.0375882
rPAD/307 PAD:14164 PAD:14167 0.0751765
rPAD/308 PAD:14161 PAD:14164 0.0375882
rPAD/309 PAD:14154 PAD:14157 0.0375882
rPAD/310 PAD:14151 PAD:14154 0.0751765
rPAD/311 PAD:14148 PAD:14151 0.0375882
rPAD/312 PAD:14145 PAD:14148 0.0751765
rPAD/313 PAD:14140 PAD:14143 0.0751765
rPAD/314 PAD:14131 PAD:14134 0.0375882
rPAD/315 PAD:14128 PAD:14131 0.0751765
rPAD/316 PAD:14125 PAD:14128 0.0375882
rPAD/317 PAD:14122 PAD:14125 0.0751765
rPAD/318 PAD:14119 PAD:14122 0.0375882
rPAD/319 PAD:14110 PAD:14113 0.0751765
rPAD/320 PAD:14107 PAD:14110 0.0375882
rPAD/321 PAD:14104 PAD:14107 0.0751765
rPAD/322 PAD:14101 PAD:14104 0.0375882
rPAD/323 PAD:14098 PAD:14101 0.0751765
rPAD/324 PAD:14095 PAD:14098 0.0375882
rPAD/325 PAD:14092 PAD:17014 0.0283817
rPAD/326 PAD:14092 PAD:14095 0.0751765
rPAD/327 PAD:14089 PAD:15121 0.0067651
rPAD/328 PAD:14089 PAD:15125 0.0381745
rPAD/329 PAD:14087 PAD:16658 0.0100588
rPAD/330 PAD:14084 PAD:14087 0.0751765
rPAD/331 PAD:14081 PAD:14084 0.0375882
rPAD/332 PAD:14072 PAD:14075 0.0751765
rPAD/333 PAD:14069 PAD:14072 0.0375882
rPAD/334 PAD:14066 PAD:14069 0.0751765
rPAD/335 PAD:14063 PAD:14066 0.0375882
rPAD/336 PAD:14060 PAD:14063 0.0751765
rPAD/337 PAD:14057 PAD:14060 0.0375882
rPAD/338 PAD:14054 PAD:14057 0.0751765
rPAD/339 PAD:14051 PAD:14054 0.0375882
rPAD/340 PAD:14048 PAD:14051 0.0751765
rPAD/341 PAD:14045 PAD:14048 0.0375882
rPAD/342 PAD:14032 PAD:14035 0.0375882
rPAD/343 PAD:14029 PAD:14032 0.0751765
rPAD/344 PAD:14020 PAD:14023 0.0375882
rPAD/345 PAD:14015 PAD:14018 0.0375882
rPAD/346 PAD:14012 PAD:14015 0.0751765
rPAD/347 PAD:14009 PAD:14012 0.0375882
rPAD/348 PAD:14006 PAD:14009 0.0751765
rPAD/349 PAD:14003 PAD:14006 0.0375882
rPAD/350 PAD:13994 PAD:13997 0.0751765
rPAD/351 PAD:13991 PAD:13994 0.0375882
rPAD/352 PAD:13984 PAD:13987 0.0375882
rPAD/353 PAD:13981 PAD:13984 0.0751765
rPAD/354 PAD:13978 PAD:13981 0.0375882
rPAD/355 PAD:13975 PAD:13978 0.0751765
rPAD/356 PAD:13970 PAD:13973 0.0751765
rPAD/357 PAD:13961 PAD:13964 0.0375882
rPAD/358 PAD:13958 PAD:13961 0.0751765
rPAD/359 PAD:13955 PAD:13958 0.0375882
rPAD/360 PAD:13952 PAD:13955 0.0751765
rPAD/361 PAD:13949 PAD:13952 0.0375882
rPAD/362 PAD:13940 PAD:13943 0.0751765
rPAD/363 PAD:13937 PAD:13940 0.0375882
rPAD/364 PAD:13934 PAD:13937 0.0751765
rPAD/365 PAD:13931 PAD:13934 0.0375882
rPAD/366 PAD:13928 PAD:13931 0.0751765
rPAD/367 PAD:13925 PAD:13928 0.0375882
rPAD/368 PAD:13922 PAD:17012 0.0283817
rPAD/369 PAD:13922 PAD:13925 0.0751765
rPAD/370 PAD:13919 PAD:15117 0.0183624
rPAD/371 PAD:13919 PAD:15121 0.041557
rPAD/372 PAD:13917 PAD:16600 0.0100588
rPAD/373 PAD:13914 PAD:13917 0.0751765
rPAD/374 PAD:13911 PAD:13914 0.0375882
rPAD/375 PAD:13902 PAD:13905 0.0751765
rPAD/376 PAD:13899 PAD:13902 0.0375882
rPAD/377 PAD:13896 PAD:13899 0.0751765
rPAD/378 PAD:13893 PAD:13896 0.0375882
rPAD/379 PAD:13890 PAD:13893 0.0751765
rPAD/380 PAD:13887 PAD:13890 0.0375882
rPAD/381 PAD:13884 PAD:13887 0.0751765
rPAD/382 PAD:13881 PAD:13884 0.0375882
rPAD/383 PAD:13878 PAD:13881 0.0751765
rPAD/384 PAD:13875 PAD:13878 0.0375882
rPAD/385 PAD:13862 PAD:13865 0.0375882
rPAD/386 PAD:13859 PAD:13862 0.0751765
rPAD/387 PAD:13850 PAD:13853 0.0375882
rPAD/388 PAD:13845 PAD:13848 0.0375882
rPAD/389 PAD:13842 PAD:13845 0.0751765
rPAD/390 PAD:13839 PAD:13842 0.0375882
rPAD/391 PAD:13836 PAD:13839 0.0751765
rPAD/392 PAD:13833 PAD:13836 0.0375882
rPAD/393 PAD:13824 PAD:13827 0.0751765
rPAD/394 PAD:13821 PAD:13824 0.0375882
rPAD/395 PAD:13814 PAD:13817 0.0375882
rPAD/396 PAD:13811 PAD:13814 0.0751765
rPAD/397 PAD:13808 PAD:13811 0.0375882
rPAD/398 PAD:13805 PAD:13808 0.0751765
rPAD/399 PAD:13800 PAD:13803 0.0751765
rPAD/400 PAD:13791 PAD:13794 0.0375882
rPAD/401 PAD:13788 PAD:13791 0.0751765
rPAD/402 PAD:13785 PAD:13788 0.0375882
rPAD/403 PAD:13782 PAD:13785 0.0751765
rPAD/404 PAD:13779 PAD:13782 0.0375882
rPAD/405 PAD:13770 PAD:13773 0.0751765
rPAD/406 PAD:13767 PAD:13770 0.0375882
rPAD/407 PAD:13764 PAD:13767 0.0751765
rPAD/408 PAD:13761 PAD:13764 0.0375882
rPAD/409 PAD:13758 PAD:13761 0.0751765
rPAD/410 PAD:13755 PAD:13758 0.0375882
rPAD/411 PAD:13752 PAD:17009 0.0283817
rPAD/412 PAD:13752 PAD:13755 0.0751765
rPAD/413 PAD:13749 PAD:15113 0.0149799
rPAD/414 PAD:13749 PAD:15117 0.0299597
rPAD/415 PAD:13747 PAD:16542 0.0100588
rPAD/416 PAD:13744 PAD:13747 0.0751765
rPAD/417 PAD:13741 PAD:13744 0.0375882
rPAD/418 PAD:13732 PAD:13735 0.0751765
rPAD/419 PAD:13729 PAD:13732 0.0375882
rPAD/420 PAD:13726 PAD:13729 0.0751765
rPAD/421 PAD:13723 PAD:13726 0.0375882
rPAD/422 PAD:13720 PAD:13723 0.0751765
rPAD/423 PAD:13717 PAD:13720 0.0375882
rPAD/424 PAD:13714 PAD:13717 0.0751765
rPAD/425 PAD:13711 PAD:13714 0.0375882
rPAD/426 PAD:13708 PAD:13711 0.0751765
rPAD/427 PAD:13705 PAD:13708 0.0375882
rPAD/428 PAD:13692 PAD:13695 0.0375882
rPAD/429 PAD:13689 PAD:13692 0.0751765
rPAD/430 PAD:13680 PAD:13683 0.0375882
rPAD/431 PAD:13675 PAD:13678 0.0375882
rPAD/432 PAD:13672 PAD:13675 0.0751765
rPAD/433 PAD:13669 PAD:13672 0.0375882
rPAD/434 PAD:13666 PAD:13669 0.0751765
rPAD/435 PAD:13663 PAD:13666 0.0375882
rPAD/436 PAD:13654 PAD:13657 0.0751765
rPAD/437 PAD:13651 PAD:13654 0.0375882
rPAD/438 PAD:13644 PAD:13647 0.0375882
rPAD/439 PAD:13641 PAD:13644 0.0751765
rPAD/440 PAD:13638 PAD:13641 0.0375882
rPAD/441 PAD:13635 PAD:13638 0.0751765
rPAD/442 PAD:13630 PAD:13633 0.0751765
rPAD/443 PAD:13621 PAD:13624 0.0375882
rPAD/444 PAD:13618 PAD:13621 0.0751765
rPAD/445 PAD:13615 PAD:13618 0.0375882
rPAD/446 PAD:13612 PAD:13615 0.0751765
rPAD/447 PAD:13609 PAD:13612 0.0375882
rPAD/448 PAD:13600 PAD:13603 0.0751765
rPAD/449 PAD:13597 PAD:13600 0.0375882
rPAD/450 PAD:13594 PAD:13597 0.0751765
rPAD/451 PAD:13591 PAD:13594 0.0375882
rPAD/452 PAD:13588 PAD:13591 0.0751765
rPAD/453 PAD:13585 PAD:13588 0.0375882
rPAD/454 PAD:13582 PAD:17007 0.0283817
rPAD/455 PAD:13582 PAD:13585 0.0751765
rPAD/456 PAD:13579 PAD:15109 0.0115973
rPAD/457 PAD:13579 PAD:15113 0.0333423
rPAD/458 PAD:13577 PAD:16484 0.0100588
rPAD/459 PAD:13574 PAD:13577 0.0751765
rPAD/460 PAD:13571 PAD:13574 0.0375882
rPAD/461 PAD:13562 PAD:13565 0.0751765
rPAD/462 PAD:13559 PAD:13562 0.0375882
rPAD/463 PAD:13556 PAD:13559 0.0751765
rPAD/464 PAD:13553 PAD:13556 0.0375882
rPAD/465 PAD:13550 PAD:13553 0.0751765
rPAD/466 PAD:13547 PAD:13550 0.0375882
rPAD/467 PAD:13544 PAD:13547 0.0751765
rPAD/468 PAD:13541 PAD:13544 0.0375882
rPAD/469 PAD:13538 PAD:13541 0.0751765
rPAD/470 PAD:13535 PAD:13538 0.0375882
rPAD/471 PAD:13522 PAD:13525 0.0375882
rPAD/472 PAD:13519 PAD:13522 0.0751765
rPAD/473 PAD:13510 PAD:13513 0.0375882
rPAD/474 PAD:13505 PAD:13508 0.0375882
rPAD/475 PAD:13502 PAD:13505 0.0751765
rPAD/476 PAD:13499 PAD:13502 0.0375882
rPAD/477 PAD:13496 PAD:13499 0.0751765
rPAD/478 PAD:13493 PAD:13496 0.0375882
rPAD/479 PAD:13484 PAD:13487 0.0751765
rPAD/480 PAD:13481 PAD:13484 0.0375882
rPAD/481 PAD:13474 PAD:13477 0.0375882
rPAD/482 PAD:13471 PAD:13474 0.0751765
rPAD/483 PAD:13468 PAD:13471 0.0375882
rPAD/484 PAD:13465 PAD:13468 0.0751765
rPAD/485 PAD:13460 PAD:13463 0.0751765
rPAD/486 PAD:13451 PAD:13454 0.0375882
rPAD/487 PAD:13448 PAD:13451 0.0751765
rPAD/488 PAD:13445 PAD:13448 0.0375882
rPAD/489 PAD:13442 PAD:13445 0.0751765
rPAD/490 PAD:13439 PAD:13442 0.0375882
rPAD/491 PAD:13430 PAD:13433 0.0751765
rPAD/492 PAD:13427 PAD:13430 0.0375882
rPAD/493 PAD:13424 PAD:13427 0.0751765
rPAD/494 PAD:13421 PAD:13424 0.0375882
rPAD/495 PAD:13418 PAD:13421 0.0751765
rPAD/496 PAD:13415 PAD:13418 0.0375882
rPAD/497 PAD:13412 PAD:17005 0.0283817
rPAD/498 PAD:13412 PAD:13415 0.0751765
rPAD/499 PAD:13409 PAD:15105 0.00821477
rPAD/500 PAD:13409 PAD:15109 0.0367248
rPAD/501 PAD:13407 PAD:16426 0.0100588
rPAD/502 PAD:13404 PAD:13407 0.0751765
rPAD/503 PAD:13401 PAD:13404 0.0375882
rPAD/504 PAD:13392 PAD:13395 0.0751765
rPAD/505 PAD:13389 PAD:13392 0.0375882
rPAD/506 PAD:13386 PAD:13389 0.0751765
rPAD/507 PAD:13383 PAD:13386 0.0375882
rPAD/508 PAD:13380 PAD:13383 0.0751765
rPAD/509 PAD:13377 PAD:13380 0.0375882
rPAD/510 PAD:13374 PAD:13377 0.0751765
rPAD/511 PAD:13371 PAD:13374 0.0375882
rPAD/512 PAD:13368 PAD:13371 0.0751765
rPAD/513 PAD:13365 PAD:13368 0.0375882
rPAD/514 PAD:13352 PAD:13355 0.0375882
rPAD/515 PAD:13349 PAD:13352 0.0751765
rPAD/516 PAD:13340 PAD:13343 0.0375882
rPAD/517 PAD:13335 PAD:13338 0.0375882
rPAD/518 PAD:13332 PAD:13335 0.0751765
rPAD/519 PAD:13329 PAD:13332 0.0375882
rPAD/520 PAD:13326 PAD:13329 0.0751765
rPAD/521 PAD:13323 PAD:13326 0.0375882
rPAD/522 PAD:13314 PAD:13317 0.0751765
rPAD/523 PAD:13311 PAD:13314 0.0375882
rPAD/524 PAD:13304 PAD:13307 0.0375882
rPAD/525 PAD:13301 PAD:13304 0.0751765
rPAD/526 PAD:13298 PAD:13301 0.0375882
rPAD/527 PAD:13295 PAD:13298 0.0751765
rPAD/528 PAD:13290 PAD:13293 0.0751765
rPAD/529 PAD:13281 PAD:13284 0.0375882
rPAD/530 PAD:13278 PAD:13281 0.0751765
rPAD/531 PAD:13275 PAD:13278 0.0375882
rPAD/532 PAD:13272 PAD:13275 0.0751765
rPAD/533 PAD:13269 PAD:13272 0.0375882
rPAD/534 PAD:13260 PAD:13263 0.0751765
rPAD/535 PAD:13257 PAD:13260 0.0375882
rPAD/536 PAD:13254 PAD:13257 0.0751765
rPAD/537 PAD:13251 PAD:13254 0.0375882
rPAD/538 PAD:13248 PAD:13251 0.0751765
rPAD/539 PAD:13245 PAD:13248 0.0375882
rPAD/540 PAD:13242 PAD:17003 0.0283817
rPAD/541 PAD:13242 PAD:13245 0.0751765
rPAD/542 PAD:13239 PAD:15101 0.0198121
rPAD/543 PAD:13239 PAD:15105 0.0401074
rPAD/544 PAD:13237 PAD:16368 0.0100588
rPAD/545 PAD:13234 PAD:13237 0.0751765
rPAD/546 PAD:13231 PAD:13234 0.0375882
rPAD/547 PAD:13222 PAD:13225 0.0751765
rPAD/548 PAD:13219 PAD:13222 0.0375882
rPAD/549 PAD:13216 PAD:13219 0.0751765
rPAD/550 PAD:13213 PAD:13216 0.0375882
rPAD/551 PAD:13210 PAD:13213 0.0751765
rPAD/552 PAD:13207 PAD:13210 0.0375882
rPAD/553 PAD:13204 PAD:13207 0.0751765
rPAD/554 PAD:13201 PAD:13204 0.0375882
rPAD/555 PAD:13198 PAD:13201 0.0751765
rPAD/556 PAD:13195 PAD:13198 0.0375882
rPAD/557 PAD:13182 PAD:13185 0.0375882
rPAD/558 PAD:13179 PAD:13182 0.0751765
rPAD/559 PAD:13170 PAD:13173 0.0375882
rPAD/560 PAD:13165 PAD:13168 0.0375882
rPAD/561 PAD:13162 PAD:13165 0.0751765
rPAD/562 PAD:13159 PAD:13162 0.0375882
rPAD/563 PAD:13156 PAD:13159 0.0751765
rPAD/564 PAD:13153 PAD:13156 0.0375882
rPAD/565 PAD:13144 PAD:13147 0.0751765
rPAD/566 PAD:13141 PAD:13144 0.0375882
rPAD/567 PAD:13134 PAD:13137 0.0375882
rPAD/568 PAD:13131 PAD:13134 0.0751765
rPAD/569 PAD:13128 PAD:13131 0.0375882
rPAD/570 PAD:13125 PAD:13128 0.0751765
rPAD/571 PAD:13120 PAD:13123 0.0751765
rPAD/572 PAD:13111 PAD:13114 0.0375882
rPAD/573 PAD:13108 PAD:13111 0.0751765
rPAD/574 PAD:13105 PAD:13108 0.0375882
rPAD/575 PAD:13102 PAD:13105 0.0751765
rPAD/576 PAD:13099 PAD:13102 0.0375882
rPAD/577 PAD:13090 PAD:13093 0.0751765
rPAD/578 PAD:13087 PAD:13090 0.0375882
rPAD/579 PAD:13084 PAD:13087 0.0751765
rPAD/580 PAD:13081 PAD:13084 0.0375882
rPAD/581 PAD:13078 PAD:13081 0.0751765
rPAD/582 PAD:13075 PAD:13078 0.0375882
rPAD/583 PAD:13072 PAD:17001 0.0283817
rPAD/584 PAD:13072 PAD:13075 0.0751765
rPAD/585 PAD:13069 PAD:15097 0.0164295
rPAD/586 PAD:13069 PAD:15101 0.0285101
rPAD/587 PAD:13067 PAD:16310 0.0100588
rPAD/588 PAD:13064 PAD:13067 0.0751765
rPAD/589 PAD:13061 PAD:13064 0.0375882
rPAD/590 PAD:13052 PAD:13055 0.0751765
rPAD/591 PAD:13049 PAD:13052 0.0375882
rPAD/592 PAD:13046 PAD:13049 0.0751765
rPAD/593 PAD:13043 PAD:13046 0.0375882
rPAD/594 PAD:13040 PAD:13043 0.0751765
rPAD/595 PAD:13037 PAD:13040 0.0375882
rPAD/596 PAD:13034 PAD:13037 0.0751765
rPAD/597 PAD:13031 PAD:13034 0.0375882
rPAD/598 PAD:13028 PAD:13031 0.0751765
rPAD/599 PAD:13025 PAD:13028 0.0375882
rPAD/600 PAD:13012 PAD:13015 0.0375882
rPAD/601 PAD:13009 PAD:13012 0.0751765
rPAD/602 PAD:13000 PAD:13003 0.0375882
rPAD/603 PAD:12995 PAD:12998 0.0375882
rPAD/604 PAD:12992 PAD:12995 0.0751765
rPAD/605 PAD:12989 PAD:12992 0.0375882
rPAD/606 PAD:12986 PAD:12989 0.0751765
rPAD/607 PAD:12983 PAD:12986 0.0375882
rPAD/608 PAD:12974 PAD:12977 0.0751765
rPAD/609 PAD:12971 PAD:12974 0.0375882
rPAD/610 PAD:12964 PAD:12967 0.0375882
rPAD/611 PAD:12961 PAD:12964 0.0751765
rPAD/612 PAD:12958 PAD:12961 0.0375882
rPAD/613 PAD:12955 PAD:12958 0.0751765
rPAD/614 PAD:12950 PAD:12953 0.0751765
rPAD/615 PAD:12941 PAD:12944 0.0375882
rPAD/616 PAD:12938 PAD:12941 0.0751765
rPAD/617 PAD:12935 PAD:12938 0.0375882
rPAD/618 PAD:12932 PAD:12935 0.0751765
rPAD/619 PAD:12929 PAD:12932 0.0375882
rPAD/620 PAD:12920 PAD:12923 0.0751765
rPAD/621 PAD:12917 PAD:12920 0.0375882
rPAD/622 PAD:12914 PAD:12917 0.0751765
rPAD/623 PAD:12911 PAD:12914 0.0375882
rPAD/624 PAD:12908 PAD:12911 0.0751765
rPAD/625 PAD:12905 PAD:12908 0.0375882
rPAD/626 PAD:12902 PAD:16999 0.0283817
rPAD/627 PAD:12902 PAD:12905 0.0751765
rPAD/628 PAD:12899 PAD:15097 0.0318926
rPAD/629 PAD:12897 PAD:16252 0.0100588
rPAD/630 PAD:12894 PAD:12897 0.0751765
rPAD/631 PAD:12891 PAD:12894 0.0375882
rPAD/632 PAD:12882 PAD:12885 0.0751765
rPAD/633 PAD:12879 PAD:12882 0.0375882
rPAD/634 PAD:12876 PAD:12879 0.0751765
rPAD/635 PAD:12873 PAD:12876 0.0375882
rPAD/636 PAD:12870 PAD:12873 0.0751765
rPAD/637 PAD:12867 PAD:12870 0.0375882
rPAD/638 PAD:12864 PAD:12867 0.0751765
rPAD/639 PAD:12861 PAD:12864 0.0375882
rPAD/640 PAD:12858 PAD:12861 0.0751765
rPAD/641 PAD:12855 PAD:12858 0.0375882
rPAD/642 PAD:12842 PAD:12845 0.0375882
rPAD/643 PAD:12839 PAD:12842 0.0751765
rPAD/644 PAD:12830 PAD:12833 0.0375882
rPAD/645 PAD:12825 PAD:12828 0.0375882
rPAD/646 PAD:12822 PAD:12825 0.0751765
rPAD/647 PAD:12819 PAD:12822 0.0375882
rPAD/648 PAD:12816 PAD:12819 0.0751765
rPAD/649 PAD:12813 PAD:12816 0.0375882
rPAD/650 PAD:12804 PAD:12807 0.0751765
rPAD/651 PAD:12801 PAD:12804 0.0375882
rPAD/652 PAD:12794 PAD:12797 0.0375882
rPAD/653 PAD:12791 PAD:12794 0.0751765
rPAD/654 PAD:12788 PAD:12791 0.0375882
rPAD/655 PAD:12785 PAD:12788 0.0751765
rPAD/656 PAD:12780 PAD:12783 0.0751765
rPAD/657 PAD:12771 PAD:12774 0.0375882
rPAD/658 PAD:12768 PAD:12771 0.0751765
rPAD/659 PAD:12765 PAD:12768 0.0375882
rPAD/660 PAD:12762 PAD:12765 0.0751765
rPAD/661 PAD:12759 PAD:12762 0.0375882
rPAD/662 PAD:12750 PAD:12753 0.0751765
rPAD/663 PAD:12747 PAD:12750 0.0375882
rPAD/664 PAD:12744 PAD:12747 0.0751765
rPAD/665 PAD:12741 PAD:12744 0.0375882
rPAD/666 PAD:12738 PAD:12741 0.0751765
rPAD/667 PAD:12735 PAD:12738 0.0375882
rPAD/668 PAD:12732 PAD:16997 0.0283817
rPAD/669 PAD:12732 PAD:12735 0.0751765
rPAD/670 PAD:12727 PAD:16194 0.0100588
rPAD/671 PAD:12724 PAD:12727 0.0751765
rPAD/672 PAD:12721 PAD:12724 0.0375882
rPAD/673 PAD:12712 PAD:12715 0.0751765
rPAD/674 PAD:12709 PAD:12712 0.0375882
rPAD/675 PAD:12706 PAD:12709 0.0751765
rPAD/676 PAD:12703 PAD:12706 0.0375882
rPAD/677 PAD:12700 PAD:12703 0.0751765
rPAD/678 PAD:12697 PAD:12700 0.0375882
rPAD/679 PAD:12694 PAD:12697 0.0751765
rPAD/680 PAD:12691 PAD:12694 0.0375882
rPAD/681 PAD:12688 PAD:12691 0.0751765
rPAD/682 PAD:12685 PAD:12688 0.0375882
rPAD/683 PAD:12672 PAD:12675 0.0375882
rPAD/684 PAD:12669 PAD:12672 0.0751765
rPAD/685 PAD:12660 PAD:12663 0.0375882
rPAD/686 PAD:12655 PAD:12658 0.0375882
rPAD/687 PAD:12652 PAD:12655 0.0751765
rPAD/688 PAD:12649 PAD:12652 0.0375882
rPAD/689 PAD:12646 PAD:12649 0.0751765
rPAD/690 PAD:12643 PAD:12646 0.0375882
rPAD/691 PAD:12634 PAD:12637 0.0751765
rPAD/692 PAD:12631 PAD:12634 0.0375882
rPAD/693 PAD:12624 PAD:12627 0.0375882
rPAD/694 PAD:12621 PAD:12624 0.0751765
rPAD/695 PAD:12618 PAD:12621 0.0375882
rPAD/696 PAD:12615 PAD:12618 0.0751765
rPAD/697 PAD:12610 PAD:12613 0.0751765
rPAD/698 PAD:12601 PAD:12604 0.0375882
rPAD/699 PAD:12598 PAD:12601 0.0751765
rPAD/700 PAD:12595 PAD:12598 0.0375882
rPAD/701 PAD:12592 PAD:12595 0.0751765
rPAD/702 PAD:12589 PAD:12592 0.0375882
rPAD/703 PAD:12580 PAD:12583 0.0751765
rPAD/704 PAD:12577 PAD:12580 0.0375882
rPAD/705 PAD:12574 PAD:12577 0.0751765
rPAD/706 PAD:12571 PAD:12574 0.0375882
rPAD/707 PAD:12568 PAD:12571 0.0751765
rPAD/708 PAD:12565 PAD:12568 0.0375882
rPAD/709 PAD:12562 PAD:16994 0.0283817
rPAD/710 PAD:12562 PAD:12565 0.0751765
rPAD/711 PAD:12557 PAD:16136 0.0100588
rPAD/712 PAD:12554 PAD:12557 0.0751765
rPAD/713 PAD:12551 PAD:12554 0.0375882
rPAD/714 PAD:12542 PAD:12545 0.0751765
rPAD/715 PAD:12539 PAD:12542 0.0375882
rPAD/716 PAD:12536 PAD:12539 0.0751765
rPAD/717 PAD:12533 PAD:12536 0.0375882
rPAD/718 PAD:12530 PAD:12533 0.0751765
rPAD/719 PAD:12527 PAD:12530 0.0375882
rPAD/720 PAD:12524 PAD:12527 0.0751765
rPAD/721 PAD:12521 PAD:12524 0.0375882
rPAD/722 PAD:12518 PAD:12521 0.0751765
rPAD/723 PAD:12515 PAD:12518 0.0375882
rPAD/724 PAD:12502 PAD:12505 0.0375882
rPAD/725 PAD:12499 PAD:12502 0.0751765
rPAD/726 PAD:12490 PAD:12493 0.0375882
rPAD/727 PAD:12485 PAD:12488 0.0375882
rPAD/728 PAD:12482 PAD:12485 0.0751765
rPAD/729 PAD:12479 PAD:12482 0.0375882
rPAD/730 PAD:12476 PAD:12479 0.0751765
rPAD/731 PAD:12473 PAD:12476 0.0375882
rPAD/732 PAD:12464 PAD:12467 0.0751765
rPAD/733 PAD:12461 PAD:12464 0.0375882
rPAD/734 PAD:12454 PAD:12457 0.0375882
rPAD/735 PAD:12451 PAD:12454 0.0751765
rPAD/736 PAD:12448 PAD:12451 0.0375882
rPAD/737 PAD:12445 PAD:12448 0.0751765
rPAD/738 PAD:12440 PAD:12443 0.0751765
rPAD/739 PAD:12431 PAD:12434 0.0375882
rPAD/740 PAD:12428 PAD:12431 0.0751765
rPAD/741 PAD:12425 PAD:12428 0.0375882
rPAD/742 PAD:12422 PAD:12425 0.0751765
rPAD/743 PAD:12419 PAD:12422 0.0375882
rPAD/744 PAD:12410 PAD:12413 0.0751765
rPAD/745 PAD:12407 PAD:12410 0.0375882
rPAD/746 PAD:12404 PAD:12407 0.0751765
rPAD/747 PAD:12401 PAD:12404 0.0375882
rPAD/748 PAD:12398 PAD:12401 0.0751765
rPAD/749 PAD:12395 PAD:12398 0.0375882
rPAD/750 PAD:12392 PAD:16992 0.0283817
rPAD/751 PAD:12392 PAD:12395 0.0751765
rPAD/752 PAD:12387 PAD:16078 0.0100588
rPAD/753 PAD:12384 PAD:12387 0.0751765
rPAD/754 PAD:12381 PAD:12384 0.0375882
rPAD/755 PAD:12372 PAD:12375 0.0751765
rPAD/756 PAD:12369 PAD:12372 0.0375882
rPAD/757 PAD:12366 PAD:12369 0.0751765
rPAD/758 PAD:12363 PAD:12366 0.0375882
rPAD/759 PAD:12360 PAD:12363 0.0751765
rPAD/760 PAD:12357 PAD:12360 0.0375882
rPAD/761 PAD:12354 PAD:12357 0.0751765
rPAD/762 PAD:12351 PAD:12354 0.0375882
rPAD/763 PAD:12348 PAD:12351 0.0751765
rPAD/764 PAD:12345 PAD:12348 0.0375882
rPAD/765 PAD:12332 PAD:12335 0.0375882
rPAD/766 PAD:12329 PAD:12332 0.0751765
rPAD/767 PAD:12320 PAD:12323 0.0375882
rPAD/768 PAD:12315 PAD:12318 0.0375882
rPAD/769 PAD:12312 PAD:12315 0.0751765
rPAD/770 PAD:12309 PAD:12312 0.0375882
rPAD/771 PAD:12306 PAD:12309 0.0751765
rPAD/772 PAD:12303 PAD:12306 0.0375882
rPAD/773 PAD:12294 PAD:12297 0.0751765
rPAD/774 PAD:12291 PAD:12294 0.0375882
rPAD/775 PAD:12284 PAD:12287 0.0375882
rPAD/776 PAD:12281 PAD:12284 0.0751765
rPAD/777 PAD:12278 PAD:12281 0.0375882
rPAD/778 PAD:12275 PAD:12278 0.0751765
rPAD/779 PAD:12270 PAD:12273 0.0751765
rPAD/780 PAD:12261 PAD:12264 0.0375882
rPAD/781 PAD:12258 PAD:12261 0.0751765
rPAD/782 PAD:12255 PAD:12258 0.0375882
rPAD/783 PAD:12252 PAD:12255 0.0751765
rPAD/784 PAD:12249 PAD:12252 0.0375882
rPAD/785 PAD:12240 PAD:12243 0.0751765
rPAD/786 PAD:12237 PAD:12240 0.0375882
rPAD/787 PAD:12234 PAD:12237 0.0751765
rPAD/788 PAD:12231 PAD:12234 0.0375882
rPAD/789 PAD:12228 PAD:12231 0.0751765
rPAD/790 PAD:12225 PAD:12228 0.0375882
rPAD/791 PAD:12222 PAD:16990 0.0283817
rPAD/792 PAD:12222 PAD:12225 0.0751765
rPAD/793 PAD:12217 PAD:16020 0.0100588
rPAD/794 PAD:12214 PAD:12217 0.0751765
rPAD/795 PAD:12211 PAD:12214 0.0375882
rPAD/796 PAD:12202 PAD:12205 0.0751765
rPAD/797 PAD:12199 PAD:12202 0.0375882
rPAD/798 PAD:12196 PAD:12199 0.0751765
rPAD/799 PAD:12193 PAD:12196 0.0375882
rPAD/800 PAD:12190 PAD:12193 0.0751765
rPAD/801 PAD:12187 PAD:12190 0.0375882
rPAD/802 PAD:12184 PAD:12187 0.0751765
rPAD/803 PAD:12181 PAD:12184 0.0375882
rPAD/804 PAD:12178 PAD:12181 0.0751765
rPAD/805 PAD:12175 PAD:12178 0.0375882
rPAD/806 PAD:12162 PAD:12165 0.0375882
rPAD/807 PAD:12159 PAD:12162 0.0751765
rPAD/808 PAD:12150 PAD:12153 0.0375882
rPAD/809 PAD:12145 PAD:12148 0.0375882
rPAD/810 PAD:12142 PAD:12145 0.0751765
rPAD/811 PAD:12139 PAD:12142 0.0375882
rPAD/812 PAD:12136 PAD:12139 0.0751765
rPAD/813 PAD:12133 PAD:12136 0.0375882
rPAD/814 PAD:12124 PAD:12127 0.0751765
rPAD/815 PAD:12121 PAD:12124 0.0375882
rPAD/816 PAD:12114 PAD:12117 0.0375882
rPAD/817 PAD:12111 PAD:12114 0.0751765
rPAD/818 PAD:12108 PAD:12111 0.0375882
rPAD/819 PAD:12105 PAD:12108 0.0751765
rPAD/820 PAD:12100 PAD:12103 0.0751765
rPAD/821 PAD:12091 PAD:12094 0.0375882
rPAD/822 PAD:12088 PAD:12091 0.0751765
rPAD/823 PAD:12085 PAD:12088 0.0375882
rPAD/824 PAD:12082 PAD:12085 0.0751765
rPAD/825 PAD:12079 PAD:12082 0.0375882
rPAD/826 PAD:12070 PAD:12073 0.0751765
rPAD/827 PAD:12067 PAD:12070 0.0375882
rPAD/828 PAD:12064 PAD:12067 0.0751765
rPAD/829 PAD:12061 PAD:12064 0.0375882
rPAD/830 PAD:12058 PAD:12061 0.0751765
rPAD/831 PAD:12055 PAD:12058 0.0375882
rPAD/832 PAD:12052 PAD:16988 0.0283817
rPAD/833 PAD:12052 PAD:12055 0.0751765
rPAD/834 PAD:12049 PAD:15073 0.0111141
rPAD/835 PAD:12047 PAD:15962 0.0100588
rPAD/836 PAD:12044 PAD:12047 0.0751765
rPAD/837 PAD:12041 PAD:12044 0.0375882
rPAD/838 PAD:12032 PAD:12035 0.0751765
rPAD/839 PAD:12029 PAD:12032 0.0375882
rPAD/840 PAD:12026 PAD:12029 0.0751765
rPAD/841 PAD:12023 PAD:12026 0.0375882
rPAD/842 PAD:12020 PAD:12023 0.0751765
rPAD/843 PAD:12017 PAD:12020 0.0375882
rPAD/844 PAD:12014 PAD:12017 0.0751765
rPAD/845 PAD:12011 PAD:12014 0.0375882
rPAD/846 PAD:12008 PAD:12011 0.0751765
rPAD/847 PAD:12005 PAD:12008 0.0375882
rPAD/848 PAD:11992 PAD:11995 0.0375882
rPAD/849 PAD:11989 PAD:11992 0.0751765
rPAD/850 PAD:11980 PAD:11983 0.0375882
rPAD/851 PAD:11975 PAD:11978 0.0375882
rPAD/852 PAD:11972 PAD:11975 0.0751765
rPAD/853 PAD:11969 PAD:11972 0.0375882
rPAD/854 PAD:11966 PAD:11969 0.0751765
rPAD/855 PAD:11963 PAD:11966 0.0375882
rPAD/856 PAD:11954 PAD:11957 0.0751765
rPAD/857 PAD:11951 PAD:11954 0.0375882
rPAD/858 PAD:11944 PAD:11947 0.0375882
rPAD/859 PAD:11941 PAD:11944 0.0751765
rPAD/860 PAD:11938 PAD:11941 0.0375882
rPAD/861 PAD:11935 PAD:11938 0.0751765
rPAD/862 PAD:11930 PAD:11933 0.0751765
rPAD/863 PAD:11921 PAD:11924 0.0375882
rPAD/864 PAD:11918 PAD:11921 0.0751765
rPAD/865 PAD:11915 PAD:11918 0.0375882
rPAD/866 PAD:11912 PAD:11915 0.0751765
rPAD/867 PAD:11909 PAD:11912 0.0375882
rPAD/868 PAD:11900 PAD:11903 0.0751765
rPAD/869 PAD:11897 PAD:11900 0.0375882
rPAD/870 PAD:11894 PAD:11897 0.0751765
rPAD/871 PAD:11891 PAD:11894 0.0375882
rPAD/872 PAD:11888 PAD:11891 0.0751765
rPAD/873 PAD:11885 PAD:11888 0.0375882
rPAD/874 PAD:11882 PAD:16986 0.0283817
rPAD/875 PAD:11882 PAD:11885 0.0751765
rPAD/876 PAD:11879 PAD:15069 0.0227114
rPAD/877 PAD:11879 PAD:15073 0.0372081
rPAD/878 PAD:11877 PAD:15904 0.0100588
rPAD/879 PAD:11874 PAD:11877 0.0751765
rPAD/880 PAD:11871 PAD:11874 0.0375882
rPAD/881 PAD:11862 PAD:11865 0.0751765
rPAD/882 PAD:11859 PAD:11862 0.0375882
rPAD/883 PAD:11856 PAD:11859 0.0751765
rPAD/884 PAD:11853 PAD:11856 0.0375882
rPAD/885 PAD:11850 PAD:11853 0.0751765
rPAD/886 PAD:11847 PAD:11850 0.0375882
rPAD/887 PAD:11844 PAD:11847 0.0751765
rPAD/888 PAD:11841 PAD:11844 0.0375882
rPAD/889 PAD:11838 PAD:11841 0.0751765
rPAD/890 PAD:11835 PAD:11838 0.0375882
rPAD/891 PAD:11822 PAD:11825 0.0375882
rPAD/892 PAD:11819 PAD:11822 0.0751765
rPAD/893 PAD:11810 PAD:11813 0.0375882
rPAD/894 PAD:11805 PAD:11808 0.0375882
rPAD/895 PAD:11802 PAD:11805 0.0751765
rPAD/896 PAD:11799 PAD:11802 0.0375882
rPAD/897 PAD:11796 PAD:11799 0.0751765
rPAD/898 PAD:11793 PAD:11796 0.0375882
rPAD/899 PAD:11784 PAD:11787 0.0751765
rPAD/900 PAD:11781 PAD:11784 0.0375882
rPAD/901 PAD:11774 PAD:11777 0.0375882
rPAD/902 PAD:11771 PAD:11774 0.0751765
rPAD/903 PAD:11768 PAD:11771 0.0375882
rPAD/904 PAD:11765 PAD:11768 0.0751765
rPAD/905 PAD:11760 PAD:11763 0.0751765
rPAD/906 PAD:11751 PAD:11754 0.0375882
rPAD/907 PAD:11748 PAD:11751 0.0751765
rPAD/908 PAD:11745 PAD:11748 0.0375882
rPAD/909 PAD:11742 PAD:11745 0.0751765
rPAD/910 PAD:11739 PAD:11742 0.0375882
rPAD/911 PAD:11730 PAD:11733 0.0751765
rPAD/912 PAD:11727 PAD:11730 0.0375882
rPAD/913 PAD:11724 PAD:11727 0.0751765
rPAD/914 PAD:11721 PAD:11724 0.0375882
rPAD/915 PAD:11718 PAD:11721 0.0751765
rPAD/916 PAD:11715 PAD:11718 0.0375882
rPAD/917 PAD:11712 PAD:16984 0.0283817
rPAD/918 PAD:11712 PAD:11715 0.0751765
rPAD/919 PAD:11709 PAD:15065 0.0193289
rPAD/920 PAD:11709 PAD:15069 0.0256107
rPAD/921 PAD:11707 PAD:15846 0.0100588
rPAD/922 PAD:11704 PAD:11707 0.0751765
rPAD/923 PAD:11701 PAD:11704 0.0375882
rPAD/924 PAD:11692 PAD:11695 0.0751765
rPAD/925 PAD:11689 PAD:11692 0.0375882
rPAD/926 PAD:11686 PAD:11689 0.0751765
rPAD/927 PAD:11683 PAD:11686 0.0375882
rPAD/928 PAD:11680 PAD:11683 0.0751765
rPAD/929 PAD:11677 PAD:11680 0.0375882
rPAD/930 PAD:11674 PAD:11677 0.0751765
rPAD/931 PAD:11671 PAD:11674 0.0375882
rPAD/932 PAD:11668 PAD:11671 0.0751765
rPAD/933 PAD:11665 PAD:11668 0.0375882
rPAD/934 PAD:11652 PAD:11655 0.0375882
rPAD/935 PAD:11649 PAD:11652 0.0751765
rPAD/936 PAD:11640 PAD:11643 0.0375882
rPAD/937 PAD:11635 PAD:11638 0.0375882
rPAD/938 PAD:11632 PAD:11635 0.0751765
rPAD/939 PAD:11629 PAD:11632 0.0375882
rPAD/940 PAD:11626 PAD:11629 0.0751765
rPAD/941 PAD:11623 PAD:11626 0.0375882
rPAD/942 PAD:11614 PAD:11617 0.0751765
rPAD/943 PAD:11611 PAD:11614 0.0375882
rPAD/944 PAD:11604 PAD:11607 0.0375882
rPAD/945 PAD:11601 PAD:11604 0.0751765
rPAD/946 PAD:11598 PAD:11601 0.0375882
rPAD/947 PAD:11595 PAD:11598 0.0751765
rPAD/948 PAD:11590 PAD:11593 0.0751765
rPAD/949 PAD:11581 PAD:11584 0.0375882
rPAD/950 PAD:11578 PAD:11581 0.0751765
rPAD/951 PAD:11575 PAD:11578 0.0375882
rPAD/952 PAD:11572 PAD:11575 0.0751765
rPAD/953 PAD:11569 PAD:11572 0.0375882
rPAD/954 PAD:11560 PAD:11563 0.0751765
rPAD/955 PAD:11557 PAD:11560 0.0375882
rPAD/956 PAD:11554 PAD:11557 0.0751765
rPAD/957 PAD:11551 PAD:11554 0.0375882
rPAD/958 PAD:11548 PAD:11551 0.0751765
rPAD/959 PAD:11545 PAD:11548 0.0375882
rPAD/960 PAD:11542 PAD:16982 0.0283817
rPAD/961 PAD:11542 PAD:11545 0.0751765
rPAD/962 PAD:11539 PAD:15061 0.0159463
rPAD/963 PAD:11539 PAD:15065 0.0289933
rPAD/964 PAD:11537 PAD:15788 0.0100588
rPAD/965 PAD:11534 PAD:11537 0.0751765
rPAD/966 PAD:11531 PAD:11534 0.0375882
rPAD/967 PAD:11522 PAD:11525 0.0751765
rPAD/968 PAD:11519 PAD:11522 0.0375882
rPAD/969 PAD:11516 PAD:11519 0.0751765
rPAD/970 PAD:11513 PAD:11516 0.0375882
rPAD/971 PAD:11510 PAD:11513 0.0751765
rPAD/972 PAD:11507 PAD:11510 0.0375882
rPAD/973 PAD:11504 PAD:11507 0.0751765
rPAD/974 PAD:11501 PAD:11504 0.0375882
rPAD/975 PAD:11498 PAD:11501 0.0751765
rPAD/976 PAD:11495 PAD:11498 0.0375882
rPAD/977 PAD:11482 PAD:11485 0.0375882
rPAD/978 PAD:11479 PAD:11482 0.0751765
rPAD/979 PAD:11470 PAD:11473 0.0375882
rPAD/980 PAD:11465 PAD:11468 0.0375882
rPAD/981 PAD:11462 PAD:11465 0.0751765
rPAD/982 PAD:11459 PAD:11462 0.0375882
rPAD/983 PAD:11456 PAD:11459 0.0751765
rPAD/984 PAD:11453 PAD:11456 0.0375882
rPAD/985 PAD:11444 PAD:11447 0.0751765
rPAD/986 PAD:11441 PAD:11444 0.0375882
rPAD/987 PAD:11434 PAD:11437 0.0375882
rPAD/988 PAD:11431 PAD:11434 0.0751765
rPAD/989 PAD:11428 PAD:11431 0.0375882
rPAD/990 PAD:11425 PAD:11428 0.0751765
rPAD/991 PAD:11420 PAD:11423 0.0751765
rPAD/992 PAD:11411 PAD:11414 0.0375882
rPAD/993 PAD:11408 PAD:11411 0.0751765
rPAD/994 PAD:11405 PAD:11408 0.0375882
rPAD/995 PAD:11402 PAD:11405 0.0751765
rPAD/996 PAD:11399 PAD:11402 0.0375882
rPAD/997 PAD:11390 PAD:11393 0.0751765
rPAD/998 PAD:11387 PAD:11390 0.0375882
rPAD/999 PAD:11384 PAD:11387 0.0751765
rPAD/1000 PAD:11381 PAD:11384 0.0375882
rPAD/1001 PAD:11378 PAD:11381 0.0751765
rPAD/1002 PAD:11375 PAD:11378 0.0375882
rPAD/1003 PAD:11372 PAD:16979 0.0283817
rPAD/1004 PAD:11372 PAD:11375 0.0751765
rPAD/1005 PAD:11369 PAD:15057 0.0125638
rPAD/1006 PAD:11369 PAD:15061 0.0323758
rPAD/1007 PAD:11367 PAD:15730 0.0100588
rPAD/1008 PAD:11364 PAD:11367 0.0751765
rPAD/1009 PAD:11361 PAD:11364 0.0375882
rPAD/1010 PAD:11352 PAD:11355 0.0751765
rPAD/1011 PAD:11349 PAD:11352 0.0375882
rPAD/1012 PAD:11346 PAD:11349 0.0751765
rPAD/1013 PAD:11343 PAD:11346 0.0375882
rPAD/1014 PAD:11340 PAD:11343 0.0751765
rPAD/1015 PAD:11337 PAD:11340 0.0375882
rPAD/1016 PAD:11334 PAD:11337 0.0751765
rPAD/1017 PAD:11331 PAD:11334 0.0375882
rPAD/1018 PAD:11328 PAD:11331 0.0751765
rPAD/1019 PAD:11325 PAD:11328 0.0375882
rPAD/1020 PAD:11312 PAD:11315 0.0375882
rPAD/1021 PAD:11309 PAD:11312 0.0751765
rPAD/1022 PAD:11300 PAD:11303 0.0375882
rPAD/1023 PAD:11295 PAD:11298 0.0375882
rPAD/1024 PAD:11292 PAD:11295 0.0751765
rPAD/1025 PAD:11289 PAD:11292 0.0375882
rPAD/1026 PAD:11286 PAD:11289 0.0751765
rPAD/1027 PAD:11283 PAD:11286 0.0375882
rPAD/1028 PAD:11274 PAD:11277 0.0751765
rPAD/1029 PAD:11271 PAD:11274 0.0375882
rPAD/1030 PAD:11264 PAD:11267 0.0375882
rPAD/1031 PAD:11261 PAD:11264 0.0751765
rPAD/1032 PAD:11258 PAD:11261 0.0375882
rPAD/1033 PAD:11255 PAD:11258 0.0751765
rPAD/1034 PAD:11250 PAD:11253 0.0751765
rPAD/1035 PAD:11241 PAD:11244 0.0375882
rPAD/1036 PAD:11238 PAD:11241 0.0751765
rPAD/1037 PAD:11235 PAD:11238 0.0375882
rPAD/1038 PAD:11232 PAD:11235 0.0751765
rPAD/1039 PAD:11229 PAD:11232 0.0375882
rPAD/1040 PAD:11220 PAD:11223 0.0751765
rPAD/1041 PAD:11217 PAD:11220 0.0375882
rPAD/1042 PAD:11214 PAD:11217 0.0751765
rPAD/1043 PAD:11211 PAD:11214 0.0375882
rPAD/1044 PAD:11208 PAD:11211 0.0751765
rPAD/1045 PAD:11205 PAD:11208 0.0375882
rPAD/1046 PAD:11202 PAD:16978 0.0283817
rPAD/1047 PAD:11202 PAD:11205 0.0751765
rPAD/1048 PAD:11199 PAD:15053 0.0241611
rPAD/1049 PAD:11199 PAD:15057 0.0357584
rPAD/1050 PAD:11197 PAD:15672 0.0100588
rPAD/1051 PAD:11194 PAD:11197 0.0751765
rPAD/1052 PAD:11191 PAD:11194 0.0375882
rPAD/1053 PAD:11182 PAD:11185 0.0751765
rPAD/1054 PAD:11179 PAD:11182 0.0375882
rPAD/1055 PAD:11176 PAD:11179 0.0751765
rPAD/1056 PAD:11173 PAD:11176 0.0375882
rPAD/1057 PAD:11170 PAD:11173 0.0751765
rPAD/1058 PAD:11167 PAD:11170 0.0375882
rPAD/1059 PAD:11164 PAD:11167 0.0751765
rPAD/1060 PAD:11161 PAD:11164 0.0375882
rPAD/1061 PAD:11158 PAD:11161 0.0751765
rPAD/1062 PAD:11155 PAD:11158 0.0375882
rPAD/1063 PAD:11142 PAD:11145 0.0375882
rPAD/1064 PAD:11139 PAD:11142 0.0751765
rPAD/1065 PAD:11130 PAD:11133 0.0375882
rPAD/1066 PAD:11125 PAD:11128 0.0375882
rPAD/1067 PAD:11122 PAD:11125 0.0751765
rPAD/1068 PAD:11119 PAD:11122 0.0375882
rPAD/1069 PAD:11116 PAD:11119 0.0751765
rPAD/1070 PAD:11113 PAD:11116 0.0375882
rPAD/1071 PAD:11104 PAD:11107 0.0751765
rPAD/1072 PAD:11101 PAD:11104 0.0375882
rPAD/1073 PAD:11094 PAD:11097 0.0375882
rPAD/1074 PAD:11091 PAD:11094 0.0751765
rPAD/1075 PAD:11088 PAD:11091 0.0375882
rPAD/1076 PAD:11085 PAD:11088 0.0751765
rPAD/1077 PAD:11080 PAD:11083 0.0751765
rPAD/1078 PAD:11071 PAD:11074 0.0375882
rPAD/1079 PAD:11068 PAD:11071 0.0751765
rPAD/1080 PAD:11065 PAD:11068 0.0375882
rPAD/1081 PAD:11062 PAD:11065 0.0751765
rPAD/1082 PAD:11059 PAD:11062 0.0375882
rPAD/1083 PAD:11050 PAD:11053 0.0751765
rPAD/1084 PAD:11047 PAD:11050 0.0375882
rPAD/1085 PAD:11044 PAD:11047 0.0751765
rPAD/1086 PAD:11041 PAD:11044 0.0375882
rPAD/1087 PAD:11038 PAD:11041 0.0751765
rPAD/1088 PAD:11035 PAD:11038 0.0375882
rPAD/1089 PAD:11032 PAD:16975 0.0283817
rPAD/1090 PAD:11032 PAD:11035 0.0751765
rPAD/1091 PAD:11029 PAD:15049 0.0207785
rPAD/1092 PAD:11029 PAD:15053 0.0241611
rPAD/1093 PAD:11027 PAD:15614 0.0100588
rPAD/1094 PAD:11024 PAD:11027 0.0751765
rPAD/1095 PAD:11021 PAD:11024 0.0375882
rPAD/1096 PAD:11012 PAD:11015 0.0751765
rPAD/1097 PAD:11009 PAD:11012 0.0375882
rPAD/1098 PAD:11006 PAD:11009 0.0751765
rPAD/1099 PAD:11003 PAD:11006 0.0375882
rPAD/1100 PAD:11000 PAD:11003 0.0751765
rPAD/1101 PAD:10997 PAD:11000 0.0375882
rPAD/1102 PAD:10994 PAD:10997 0.0751765
rPAD/1103 PAD:10991 PAD:10994 0.0375882
rPAD/1104 PAD:10988 PAD:10991 0.0751765
rPAD/1105 PAD:10985 PAD:10988 0.0375882
rPAD/1106 PAD:10972 PAD:10975 0.0375882
rPAD/1107 PAD:10969 PAD:10972 0.0751765
rPAD/1108 PAD:10960 PAD:10963 0.0375882
rPAD/1109 PAD:10955 PAD:10958 0.0375882
rPAD/1110 PAD:10952 PAD:10955 0.0751765
rPAD/1111 PAD:10949 PAD:10952 0.0375882
rPAD/1112 PAD:10946 PAD:10949 0.0751765
rPAD/1113 PAD:10943 PAD:10946 0.0375882
rPAD/1114 PAD:10934 PAD:10937 0.0751765
rPAD/1115 PAD:10931 PAD:10934 0.0375882
rPAD/1116 PAD:10924 PAD:10927 0.0375882
rPAD/1117 PAD:10921 PAD:10924 0.0751765
rPAD/1118 PAD:10918 PAD:10921 0.0375882
rPAD/1119 PAD:10915 PAD:10918 0.0751765
rPAD/1120 PAD:10910 PAD:10913 0.0751765
rPAD/1121 PAD:10901 PAD:10904 0.0375882
rPAD/1122 PAD:10898 PAD:10901 0.0751765
rPAD/1123 PAD:10895 PAD:10898 0.0375882
rPAD/1124 PAD:10892 PAD:10895 0.0751765
rPAD/1125 PAD:10889 PAD:10892 0.0375882
rPAD/1126 PAD:10880 PAD:10883 0.0751765
rPAD/1127 PAD:10877 PAD:10880 0.0375882
rPAD/1128 PAD:10874 PAD:10877 0.0751765
rPAD/1129 PAD:10871 PAD:10874 0.0375882
rPAD/1130 PAD:10868 PAD:10871 0.0751765
rPAD/1131 PAD:10865 PAD:10868 0.0375882
rPAD/1132 PAD:10862 PAD:16973 0.0283817
rPAD/1133 PAD:10862 PAD:10865 0.0751765
rPAD/1134 PAD:10859 PAD:15045 0.017396
rPAD/1135 PAD:10859 PAD:15049 0.0275436
rPAD/1136 PAD:10857 PAD:15556 0.0100588
rPAD/1137 PAD:10854 PAD:10857 0.0751765
rPAD/1138 PAD:10851 PAD:10854 0.0375882
rPAD/1139 PAD:10842 PAD:10845 0.0751765
rPAD/1140 PAD:10839 PAD:10842 0.0375882
rPAD/1141 PAD:10836 PAD:10839 0.0751765
rPAD/1142 PAD:10833 PAD:10836 0.0375882
rPAD/1143 PAD:10830 PAD:10833 0.0751765
rPAD/1144 PAD:10827 PAD:10830 0.0375882
rPAD/1145 PAD:10824 PAD:10827 0.0751765
rPAD/1146 PAD:10821 PAD:10824 0.0375882
rPAD/1147 PAD:10818 PAD:10821 0.0751765
rPAD/1148 PAD:10815 PAD:10818 0.0375882
rPAD/1149 PAD:10802 PAD:10805 0.0375882
rPAD/1150 PAD:10799 PAD:10802 0.0751765
rPAD/1151 PAD:10790 PAD:10793 0.0375882
rPAD/1152 PAD:10785 PAD:10788 0.0375882
rPAD/1153 PAD:10782 PAD:10785 0.0751765
rPAD/1154 PAD:10779 PAD:10782 0.0375882
rPAD/1155 PAD:10776 PAD:10779 0.0751765
rPAD/1156 PAD:10773 PAD:10776 0.0375882
rPAD/1157 PAD:10764 PAD:10767 0.0751765
rPAD/1158 PAD:10761 PAD:10764 0.0375882
rPAD/1159 PAD:10754 PAD:10757 0.0375882
rPAD/1160 PAD:10751 PAD:10754 0.0751765
rPAD/1161 PAD:10748 PAD:10751 0.0375882
rPAD/1162 PAD:10745 PAD:10748 0.0751765
rPAD/1163 PAD:10740 PAD:10743 0.0751765
rPAD/1164 PAD:10731 PAD:10734 0.0375882
rPAD/1165 PAD:10728 PAD:10731 0.0751765
rPAD/1166 PAD:10725 PAD:10728 0.0375882
rPAD/1167 PAD:10722 PAD:10725 0.0751765
rPAD/1168 PAD:10719 PAD:10722 0.0375882
rPAD/1169 PAD:10710 PAD:10713 0.0751765
rPAD/1170 PAD:10707 PAD:10710 0.0375882
rPAD/1171 PAD:10704 PAD:10707 0.0751765
rPAD/1172 PAD:10701 PAD:10704 0.0375882
rPAD/1173 PAD:10698 PAD:10701 0.0751765
rPAD/1174 PAD:10695 PAD:10698 0.0375882
rPAD/1175 PAD:10692 PAD:16971 0.0283817
rPAD/1176 PAD:10692 PAD:10695 0.0751765
rPAD/1177 PAD:10689 PAD:15045 0.0309262
rPAD/1178 PAD:10687 PAD:15498 0.0100588
rPAD/1179 PAD:10684 PAD:10687 0.0751765
rPAD/1180 PAD:10681 PAD:10684 0.0375882
rPAD/1181 PAD:10672 PAD:10675 0.0751765
rPAD/1182 PAD:10669 PAD:10672 0.0375882
rPAD/1183 PAD:10666 PAD:10669 0.0751765
rPAD/1184 PAD:10663 PAD:10666 0.0375882
rPAD/1185 PAD:10660 PAD:10663 0.0751765
rPAD/1186 PAD:10657 PAD:10660 0.0375882
rPAD/1187 PAD:10654 PAD:10657 0.0751765
rPAD/1188 PAD:10651 PAD:10654 0.0375882
rPAD/1189 PAD:10648 PAD:10651 0.0751765
rPAD/1190 PAD:10645 PAD:10648 0.0375882
rPAD/1191 PAD:10632 PAD:10635 0.0375882
rPAD/1192 PAD:10629 PAD:10632 0.0751765
rPAD/1193 PAD:10620 PAD:10623 0.0375882
rPAD/1194 PAD:10615 PAD:10618 0.0375882
rPAD/1195 PAD:10612 PAD:10615 0.0751765
rPAD/1196 PAD:10609 PAD:10612 0.0375882
rPAD/1197 PAD:10606 PAD:10609 0.0751765
rPAD/1198 PAD:10603 PAD:10606 0.0375882
rPAD/1199 PAD:10594 PAD:10597 0.0751765
rPAD/1200 PAD:10591 PAD:10594 0.0375882
rPAD/1201 PAD:10584 PAD:10587 0.0375882
rPAD/1202 PAD:10581 PAD:10584 0.0751765
rPAD/1203 PAD:10578 PAD:10581 0.0375882
rPAD/1204 PAD:10575 PAD:10578 0.0751765
rPAD/1205 PAD:10570 PAD:10573 0.0751765
rPAD/1206 PAD:10561 PAD:10564 0.0375882
rPAD/1207 PAD:10558 PAD:10561 0.0751765
rPAD/1208 PAD:10555 PAD:10558 0.0375882
rPAD/1209 PAD:10552 PAD:10555 0.0751765
rPAD/1210 PAD:10549 PAD:10552 0.0375882
rPAD/1211 PAD:10540 PAD:10543 0.0751765
rPAD/1212 PAD:10537 PAD:10540 0.0375882
rPAD/1213 PAD:10534 PAD:10537 0.0751765
rPAD/1214 PAD:10531 PAD:10534 0.0375882
rPAD/1215 PAD:10528 PAD:10531 0.0751765
rPAD/1216 PAD:10525 PAD:10528 0.0375882
rPAD/1217 PAD:10522 PAD:16969 0.0283817
rPAD/1218 PAD:10522 PAD:10525 0.0751765
rPAD/1219 PAD:10517 PAD:15440 0.0100588
rPAD/1220 PAD:10514 PAD:10517 0.0751765
rPAD/1221 PAD:10511 PAD:10514 0.0375882
rPAD/1222 PAD:10502 PAD:10505 0.0751765
rPAD/1223 PAD:10499 PAD:10502 0.0375882
rPAD/1224 PAD:10496 PAD:10499 0.0751765
rPAD/1225 PAD:10493 PAD:10496 0.0375882
rPAD/1226 PAD:10490 PAD:10493 0.0751765
rPAD/1227 PAD:10487 PAD:10490 0.0375882
rPAD/1228 PAD:10484 PAD:10487 0.0751765
rPAD/1229 PAD:10481 PAD:10484 0.0375882
rPAD/1230 PAD:10478 PAD:10481 0.0751765
rPAD/1231 PAD:10475 PAD:10478 0.0375882
rPAD/1232 PAD:10462 PAD:10465 0.0375882
rPAD/1233 PAD:10459 PAD:10462 0.0751765
rPAD/1234 PAD:10450 PAD:10453 0.0375882
rPAD/1235 PAD:10445 PAD:10448 0.0375882
rPAD/1236 PAD:10442 PAD:10445 0.0751765
rPAD/1237 PAD:10439 PAD:10442 0.0375882
rPAD/1238 PAD:10436 PAD:10439 0.0751765
rPAD/1239 PAD:10433 PAD:10436 0.0375882
rPAD/1240 PAD:10424 PAD:10427 0.0751765
rPAD/1241 PAD:10421 PAD:10424 0.0375882
rPAD/1242 PAD:10414 PAD:10417 0.0375882
rPAD/1243 PAD:10411 PAD:10414 0.0751765
rPAD/1244 PAD:10408 PAD:10411 0.0375882
rPAD/1245 PAD:10405 PAD:10408 0.0751765
rPAD/1246 PAD:10400 PAD:10403 0.0751765
rPAD/1247 PAD:10391 PAD:10394 0.0375882
rPAD/1248 PAD:10388 PAD:10391 0.0751765
rPAD/1249 PAD:10385 PAD:10388 0.0375882
rPAD/1250 PAD:10382 PAD:10385 0.0751765
rPAD/1251 PAD:10379 PAD:10382 0.0375882
rPAD/1252 PAD:10370 PAD:10373 0.0751765
rPAD/1253 PAD:10367 PAD:10370 0.0375882
rPAD/1254 PAD:10364 PAD:10367 0.0751765
rPAD/1255 PAD:10361 PAD:10364 0.0375882
rPAD/1256 PAD:10358 PAD:10361 0.0751765
rPAD/1257 PAD:10355 PAD:10358 0.0375882
rPAD/1258 PAD:10352 PAD:16967 0.0283817
rPAD/1259 PAD:10352 PAD:10355 0.0751765
rPAD/1260 PAD:10347 PAD:15382 0.0100588
rPAD/1261 PAD:10344 PAD:10347 0.0751765
rPAD/1262 PAD:10341 PAD:10344 0.0375882
rPAD/1263 PAD:10332 PAD:10335 0.0751765
rPAD/1264 PAD:10329 PAD:10332 0.0375882
rPAD/1265 PAD:10326 PAD:10329 0.0751765
rPAD/1266 PAD:10323 PAD:10326 0.0375882
rPAD/1267 PAD:10320 PAD:10323 0.0751765
rPAD/1268 PAD:10317 PAD:10320 0.0375882
rPAD/1269 PAD:10314 PAD:10317 0.0751765
rPAD/1270 PAD:10311 PAD:10314 0.0375882
rPAD/1271 PAD:10308 PAD:10311 0.0751765
rPAD/1272 PAD:10305 PAD:10308 0.0375882
rPAD/1273 PAD:10292 PAD:10295 0.0375882
rPAD/1274 PAD:10289 PAD:10292 0.0751765
rPAD/1275 PAD:10280 PAD:10283 0.0375882
rPAD/1276 PAD:10275 PAD:10278 0.0375882
rPAD/1277 PAD:10272 PAD:10275 0.0751765
rPAD/1278 PAD:10269 PAD:10272 0.0375882
rPAD/1279 PAD:10266 PAD:10269 0.0751765
rPAD/1280 PAD:10263 PAD:10266 0.0375882
rPAD/1281 PAD:10254 PAD:10257 0.0751765
rPAD/1282 PAD:10251 PAD:10254 0.0375882
rPAD/1283 PAD:10244 PAD:10247 0.0375882
rPAD/1284 PAD:10241 PAD:10244 0.0751765
rPAD/1285 PAD:10238 PAD:10241 0.0375882
rPAD/1286 PAD:10235 PAD:10238 0.0751765
rPAD/1287 PAD:10230 PAD:10233 0.0751765
rPAD/1288 PAD:10221 PAD:10224 0.0375882
rPAD/1289 PAD:10218 PAD:10221 0.0751765
rPAD/1290 PAD:10215 PAD:10218 0.0375882
rPAD/1291 PAD:10212 PAD:10215 0.0751765
rPAD/1292 PAD:10209 PAD:10212 0.0375882
rPAD/1293 PAD:10200 PAD:10203 0.0751765
rPAD/1294 PAD:10197 PAD:10200 0.0375882
rPAD/1295 PAD:10194 PAD:10197 0.0751765
rPAD/1296 PAD:10191 PAD:10194 0.0375882
rPAD/1297 PAD:10188 PAD:10191 0.0751765
rPAD/1298 PAD:10185 PAD:10188 0.0375882
rPAD/1299 PAD:10182 PAD:16965 0.0283817
rPAD/1300 PAD:10182 PAD:10185 0.0751765
rPAD/1301 PAD:10177 PAD:15324 0.0100588
rPAD/1302 PAD:10174 PAD:10177 0.0751765
rPAD/1303 PAD:10171 PAD:10174 0.0375882
rPAD/1304 PAD:10162 PAD:10165 0.0751765
rPAD/1305 PAD:10159 PAD:10162 0.0375882
rPAD/1306 PAD:10156 PAD:10159 0.0751765
rPAD/1307 PAD:10153 PAD:10156 0.0375882
rPAD/1308 PAD:10150 PAD:10153 0.0751765
rPAD/1309 PAD:10147 PAD:10150 0.0375882
rPAD/1310 PAD:10144 PAD:10147 0.0751765
rPAD/1311 PAD:10141 PAD:10144 0.0375882
rPAD/1312 PAD:10138 PAD:10141 0.0751765
rPAD/1313 PAD:10135 PAD:10138 0.0375882
rPAD/1314 PAD:10122 PAD:10125 0.0375882
rPAD/1315 PAD:10119 PAD:10122 0.0751765
rPAD/1316 PAD:10110 PAD:10113 0.0375882
rPAD/1317 PAD:10105 PAD:10108 0.0375882
rPAD/1318 PAD:10102 PAD:10105 0.0751765
rPAD/1319 PAD:10099 PAD:10102 0.0375882
rPAD/1320 PAD:10096 PAD:10099 0.0751765
rPAD/1321 PAD:10093 PAD:10096 0.0375882
rPAD/1322 PAD:10084 PAD:10087 0.0751765
rPAD/1323 PAD:10081 PAD:10084 0.0375882
rPAD/1324 PAD:10074 PAD:10077 0.0375882
rPAD/1325 PAD:10071 PAD:10074 0.0751765
rPAD/1326 PAD:10068 PAD:10071 0.0375882
rPAD/1327 PAD:10065 PAD:10068 0.0751765
rPAD/1328 PAD:10060 PAD:10063 0.0751765
rPAD/1329 PAD:10051 PAD:10054 0.0375882
rPAD/1330 PAD:10048 PAD:10051 0.0751765
rPAD/1331 PAD:10045 PAD:10048 0.0375882
rPAD/1332 PAD:10042 PAD:10045 0.0751765
rPAD/1333 PAD:10039 PAD:10042 0.0375882
rPAD/1334 PAD:10030 PAD:10033 0.0751765
rPAD/1335 PAD:10027 PAD:10030 0.0375882
rPAD/1336 PAD:10024 PAD:10027 0.0751765
rPAD/1337 PAD:10021 PAD:10024 0.0375882
rPAD/1338 PAD:10018 PAD:10021 0.0751765
rPAD/1339 PAD:10015 PAD:10018 0.0375882
rPAD/1340 PAD:10012 PAD:16963 0.0283817
rPAD/1341 PAD:10012 PAD:10015 0.0751765
rPAD/1342 PAD:10007 PAD:15266 0.0100588
rPAD/1343 PAD:10004 PAD:10007 0.0751765
rPAD/1344 PAD:10001 PAD:10004 0.0375882
rPAD/1345 PAD:9992 PAD:9995 0.0751765
rPAD/1346 PAD:9989 PAD:9992 0.0375882
rPAD/1347 PAD:9986 PAD:9989 0.0751765
rPAD/1348 PAD:9983 PAD:9986 0.0375882
rPAD/1349 PAD:9980 PAD:9983 0.0751765
rPAD/1350 PAD:9977 PAD:9980 0.0375882
rPAD/1351 PAD:9974 PAD:9977 0.0751765
rPAD/1352 PAD:9971 PAD:9974 0.0375882
rPAD/1353 PAD:9968 PAD:9971 0.0751765
rPAD/1354 PAD:9965 PAD:9968 0.0375882
rPAD/1355 PAD:9952 PAD:9955 0.0375882
rPAD/1356 PAD:9949 PAD:9952 0.0751765
rPAD/1357 PAD:9940 PAD:9943 0.0375882
rPAD/1358 PAD:9935 PAD:9938 0.0375882
rPAD/1359 PAD:9932 PAD:9935 0.0751765
rPAD/1360 PAD:9929 PAD:9932 0.0375882
rPAD/1361 PAD:9926 PAD:9929 0.0751765
rPAD/1362 PAD:9923 PAD:9926 0.0375882
rPAD/1363 PAD:9914 PAD:9917 0.0751765
rPAD/1364 PAD:9911 PAD:9914 0.0375882
rPAD/1365 PAD:9904 PAD:9907 0.0375882
rPAD/1366 PAD:9901 PAD:9904 0.0751765
rPAD/1367 PAD:9898 PAD:9901 0.0375882
rPAD/1368 PAD:9895 PAD:9898 0.0751765
rPAD/1369 PAD:9890 PAD:9893 0.0751765
rPAD/1370 PAD:9881 PAD:9884 0.0375882
rPAD/1371 PAD:9878 PAD:9881 0.0751765
rPAD/1372 PAD:9875 PAD:9878 0.0375882
rPAD/1373 PAD:9872 PAD:9875 0.0751765
rPAD/1374 PAD:9869 PAD:9872 0.0375882
rPAD/1375 PAD:9860 PAD:9863 0.0751765
rPAD/1376 PAD:9857 PAD:9860 0.0375882
rPAD/1377 PAD:9854 PAD:9857 0.0751765
rPAD/1378 PAD:9851 PAD:9854 0.0375882
rPAD/1379 PAD:9848 PAD:9851 0.0751765
rPAD/1380 PAD:9845 PAD:9848 0.0375882
rPAD/1381 PAD:9842 PAD:16960 0.0283817
rPAD/1382 PAD:9842 PAD:9845 0.0751765
rPAD/1383 PAD:9839 PAD:15021 0.0270604
rPAD/1384 PAD:9837 PAD:15208 0.0100588
rPAD/1385 PAD:9834 PAD:9837 0.0751765
rPAD/1386 PAD:9831 PAD:9834 0.0375882
rPAD/1387 PAD:9822 PAD:9825 0.0751765
rPAD/1388 PAD:9819 PAD:9822 0.0375882
rPAD/1389 PAD:9816 PAD:9819 0.0751765
rPAD/1390 PAD:9813 PAD:9816 0.0375882
rPAD/1391 PAD:9810 PAD:9813 0.0751765
rPAD/1392 PAD:9807 PAD:9810 0.0375882
rPAD/1393 PAD:9804 PAD:9807 0.0751765
rPAD/1394 PAD:9801 PAD:9804 0.0375882
rPAD/1395 PAD:9798 PAD:9801 0.0751765
rPAD/1396 PAD:9795 PAD:9798 0.0375882
rPAD/1397 PAD:9782 PAD:9785 0.0375882
rPAD/1398 PAD:9779 PAD:9782 0.0751765
rPAD/1399 PAD:9770 PAD:9773 0.0375882
rPAD/1400 PAD:9765 PAD:9768 0.0375882
rPAD/1401 PAD:9762 PAD:9765 0.0751765
rPAD/1402 PAD:9759 PAD:9762 0.0375882
rPAD/1403 PAD:9756 PAD:9759 0.0751765
rPAD/1404 PAD:9753 PAD:9756 0.0375882
rPAD/1405 PAD:9744 PAD:9747 0.0751765
rPAD/1406 PAD:9741 PAD:9744 0.0375882
rPAD/1407 PAD:9734 PAD:9737 0.0375882
rPAD/1408 PAD:9731 PAD:9734 0.0751765
rPAD/1409 PAD:9728 PAD:9731 0.0375882
rPAD/1410 PAD:9725 PAD:9728 0.0751765
rPAD/1411 PAD:9720 PAD:9723 0.0751765
rPAD/1412 PAD:9711 PAD:9714 0.0375882
rPAD/1413 PAD:9708 PAD:9711 0.0751765
rPAD/1414 PAD:9705 PAD:9708 0.0375882
rPAD/1415 PAD:9702 PAD:9705 0.0751765
rPAD/1416 PAD:9699 PAD:9702 0.0375882
rPAD/1417 PAD:9690 PAD:9693 0.0751765
rPAD/1418 PAD:9687 PAD:9690 0.0375882
rPAD/1419 PAD:9684 PAD:9687 0.0751765
rPAD/1420 PAD:9681 PAD:9684 0.0375882
rPAD/1421 PAD:9678 PAD:9681 0.0751765
rPAD/1422 PAD:9675 PAD:9678 0.0375882
rPAD/1423 PAD:9672 PAD:16958 0.0283817
rPAD/1424 PAD:9672 PAD:9675 0.0751765
rPAD/1425 PAD:9669 PAD:15017 0.0236779
rPAD/1426 PAD:9669 PAD:15021 0.0212617
rPAD/1427 PAD:9666 PAD:15145 0.026775
rPAD/1428 PAD:9663 PAD:9666 0.0279
rPAD/1429 PAD:9655 PAD:9658 0.01395
rPAD/1430 PAD:9644 PAD:9647 0.01395
rPAD/1431 PAD:9644 PAD:9645 0.586956
rPAD/1432 PAD:9637 PAD:9640 0.01395
rPAD/1433 PAD:9637 PAD:9638 0.586956
rPAD/1434 PAD:9634 PAD:9637 0.01395
rPAD/1435 PAD:9630 PAD:9631 0.586956
rPAD/1436 PAD:9623 PAD:9626 0.01395
rPAD/1437 PAD:9616 PAD:9619 0.01395
rPAD/1438 PAD:9616 PAD:9617 0.586956
rPAD/1439 PAD:9613 PAD:9617 0.0279
rPAD/1440 PAD:9612 PAD:9613 0.586956
rPAD/1441 PAD:9610 PAD:9613 0.01395
rPAD/1442 PAD:9606 PAD:9610 0.0279
rPAD/1443 PAD:9605 PAD:9606 0.586956
rPAD/1444 PAD:9603 PAD:9606 0.01395
rPAD/1445 PAD:9602 PAD:9605 0.01395
rPAD/1446 PAD:9602 PAD:9603 0.586956
rPAD/1447 PAD:9599 PAD:9603 0.0279
rPAD/1448 PAD:9598 PAD:9599 0.586956
rPAD/1449 PAD:9591 PAD:9594 0.01395
rPAD/1450 PAD:9587 PAD:9588 0.586956
rPAD/1451 PAD:9584 PAD:9587 0.01395
rPAD/1452 PAD:9581 PAD:9584 0.01395
rPAD/1453 PAD:9573 PAD:9574 0.586956
rPAD/1454 PAD:9570 PAD:9573 0.01395
rPAD/1455 PAD:9563 PAD:9566 0.01395
rPAD/1456 PAD:9563 PAD:9564 0.586956
rPAD/1457 PAD:9549 PAD:9552 0.01395
rPAD/1458 PAD:9545 PAD:9546 0.586956
rPAD/1459 PAD:9542 PAD:9546 0.0279
rPAD/1460 PAD:9541 PAD:9542 0.586956
rPAD/1461 PAD:9538 PAD:9541 0.01395
rPAD/1462 PAD:9534 PAD:9535 0.586956
rPAD/1463 PAD:9531 PAD:9534 0.01395
rPAD/1464 PAD:9528 PAD:9531 0.01395
rPAD/1465 PAD:9524 PAD:9525 0.586956
rPAD/1466 PAD:9517 PAD:9520 0.01395
rPAD/1467 PAD:9510 PAD:9513 0.01395
rPAD/1468 PAD:9510 PAD:9511 0.586956
rPAD/1469 PAD:9499 PAD:9500 0.586956
rPAD/1470 PAD:9496 PAD:9499 0.01395
rPAD/1471 PAD:9485 PAD:9488 0.01395
rPAD/1472 PAD:9485 PAD:9486 0.586956
rPAD/1473 PAD:9478 PAD:9481 0.01395
rPAD/1474 PAD:9475 PAD:9478 0.01395
rPAD/1475 PAD:9475 PAD:9476 0.586956
rPAD/1476 PAD:9472 PAD:9476 0.0279
rPAD/1477 PAD:9471 PAD:9472 0.586956
rPAD/1478 PAD:9464 PAD:9467 0.01395
rPAD/1479 PAD:9464 PAD:9465 0.586956
rPAD/1480 PAD:9457 PAD:9460 0.01395
rPAD/1481 PAD:9457 PAD:9458 0.586956
rPAD/1482 PAD:9454 PAD:15144 0.01035
rPAD/1483 PAD:9454 PAD:9458 0.0279
rPAD/1484 PAD:9453 PAD:9454 0.586956
rPAD/1485 PAD:9451 PAD:15008 0.0123221
rPAD/1486 PAD:9450 PAD:14822 0.00196507
rPAD/1487 PAD:9450 PAD:9453 0.01035
rPAD/1488 PAD:9449 PAD:15142 1.5
rPAD/1489 PAD:9445 PAD:14599 0.000724832
rPAD/1490 PAD:9445 PAD:15137 0.346154
rPAD/1491 PAD:9444 PAD:9445 0.346154
rPAD/1492 PAD:9442 PAD:14429 0.0314094
rPAD/1493 PAD:9442 PAD:9445 0.0599195
rPAD/1494 PAD:9442 PAD:15134 0.346154
rPAD/1495 PAD:9441 PAD:9444 0.0649971
rPAD/1496 PAD:9441 PAD:9442 0.346154
rPAD/1497 PAD:9439 PAD:9441 0.0340711
rPAD/1498 PAD:9437 PAD:9439 0.0146768
rPAD/1499 PAD:9437 PAD:15129 0.346154
rPAD/1500 PAD:9435 PAD:9437 0.0377402
rPAD/1501 PAD:9433 PAD:9435 0.0110076
rPAD/1502 PAD:9433 PAD:15125 0.346154
rPAD/1503 PAD:9431 PAD:9433 0.0414094
rPAD/1504 PAD:9429 PAD:9431 0.00733838
rPAD/1505 PAD:9429 PAD:15121 0.346154
rPAD/1506 PAD:9427 PAD:9429 0.0450786
rPAD/1507 PAD:9425 PAD:9427 0.0199185
rPAD/1508 PAD:9425 PAD:15117 0.346154
rPAD/1509 PAD:9423 PAD:9425 0.0141526
rPAD/1510 PAD:9422 PAD:9423 0.018346
rPAD/1511 PAD:9420 PAD:9422 0.0162493
rPAD/1512 PAD:9420 PAD:15113 0.346154
rPAD/1513 PAD:9418 PAD:9420 0.0361677
rPAD/1514 PAD:9416 PAD:9418 0.0125801
rPAD/1515 PAD:9416 PAD:15109 0.346154
rPAD/1516 PAD:9414 PAD:9416 0.0398369
rPAD/1517 PAD:9412 PAD:9414 0.00891089
rPAD/1518 PAD:9412 PAD:15105 0.346154
rPAD/1519 PAD:9410 PAD:9412 0.0167734
rPAD/1520 PAD:9409 PAD:9410 0.0267327
rPAD/1521 PAD:9407 PAD:9409 0.021491
rPAD/1522 PAD:9407 PAD:15101 0.346154
rPAD/1523 PAD:9405 PAD:9407 0.030926
rPAD/1524 PAD:9403 PAD:9405 0.0178218
rPAD/1525 PAD:9403 PAD:15097 0.346154
rPAD/1526 PAD:9401 PAD:9403 0.0345952
rPAD/1527 PAD:9400 PAD:12729 0.0352752
rPAD/1528 PAD:9400 PAD:12899 0.013047
rPAD/1529 PAD:9399 PAD:9401 0.0141526
rPAD/1530 PAD:9399 PAD:9400 0.346154
rPAD/1531 PAD:9397 PAD:9399 0.00314502
rPAD/1532 PAD:9396 PAD:9397 0.0351194
rPAD/1533 PAD:9395 PAD:12559 0.0386577
rPAD/1534 PAD:9395 PAD:12729 0.00966443
rPAD/1535 PAD:9395 PAD:15090 0.346154
rPAD/1536 PAD:9394 PAD:9396 0.0104834
rPAD/1537 PAD:9394 PAD:9395 0.346154
rPAD/1538 PAD:9392 PAD:9394 0.0419336
rPAD/1539 PAD:9391 PAD:12389 0.0270604
rPAD/1540 PAD:9391 PAD:12559 0.0212617
rPAD/1541 PAD:9391 PAD:15086 0.346154
rPAD/1542 PAD:9390 PAD:9392 0.0230635
rPAD/1543 PAD:9390 PAD:9391 0.346154
rPAD/1544 PAD:9388 PAD:9390 0.0293535
rPAD/1545 PAD:9387 PAD:9388 0.00891089
rPAD/1546 PAD:9386 PAD:12219 0.030443
rPAD/1547 PAD:9386 PAD:12389 0.0178792
rPAD/1548 PAD:9386 PAD:15082 0.346154
rPAD/1549 PAD:9385 PAD:9387 0.0104834
rPAD/1550 PAD:9385 PAD:9386 0.346154
rPAD/1551 PAD:9383 PAD:9385 0.0330227
rPAD/1552 PAD:9382 PAD:12049 0.0338255
rPAD/1553 PAD:9382 PAD:12219 0.0144966
rPAD/1554 PAD:9381 PAD:9383 0.0157251
rPAD/1555 PAD:9381 PAD:9382 0.346154
rPAD/1556 PAD:9379 PAD:9381 0.0366919
rPAD/1557 PAD:9377 PAD:9379 0.0120559
rPAD/1558 PAD:9377 PAD:15073 0.346154
rPAD/1559 PAD:9375 PAD:9377 0.0403611
rPAD/1560 PAD:9373 PAD:9375 0.024636
rPAD/1561 PAD:9373 PAD:15069 0.346154
rPAD/1562 PAD:9371 PAD:9373 0.027781
rPAD/1563 PAD:9370 PAD:9371 0.00104834
rPAD/1564 PAD:9368 PAD:9370 0.0199185
rPAD/1565 PAD:9368 PAD:15065 0.346154
rPAD/1566 PAD:9366 PAD:9368 0.0314502
rPAD/1567 PAD:9364 PAD:9366 0.0172976
rPAD/1568 PAD:9364 PAD:15061 0.346154
rPAD/1569 PAD:9362 PAD:9364 0.0351194
rPAD/1570 PAD:9360 PAD:9362 0.0136284
rPAD/1571 PAD:9360 PAD:15057 0.346154
rPAD/1572 PAD:9358 PAD:9360 0.0314502
rPAD/1573 PAD:9357 PAD:9358 0.00733838
rPAD/1574 PAD:9355 PAD:9357 0.0262085
rPAD/1575 PAD:9355 PAD:15053 0.346154
rPAD/1576 PAD:9353 PAD:9355 0.0262085
rPAD/1577 PAD:9351 PAD:9353 0.0225393
rPAD/1578 PAD:9351 PAD:15049 0.346154
rPAD/1579 PAD:9349 PAD:9351 0.0298777
rPAD/1580 PAD:9347 PAD:9349 0.0188701
rPAD/1581 PAD:9347 PAD:15045 0.346154
rPAD/1582 PAD:9345 PAD:9347 0.0178218
rPAD/1583 PAD:9344 PAD:9345 0.0157251
rPAD/1584 PAD:9343 PAD:10519 0.0343087
rPAD/1585 PAD:9343 PAD:10689 0.0140134
rPAD/1586 PAD:9342 PAD:9344 0.0152009
rPAD/1587 PAD:9342 PAD:9343 0.346154
rPAD/1588 PAD:9340 PAD:9342 0.0372161
rPAD/1589 PAD:9339 PAD:10349 0.0227114
rPAD/1590 PAD:9339 PAD:10519 0.0256107
rPAD/1591 PAD:9339 PAD:15038 0.346154
rPAD/1592 PAD:9338 PAD:9340 0.027781
rPAD/1593 PAD:9338 PAD:9339 0.346154
rPAD/1594 PAD:9336 PAD:9338 0.024636
rPAD/1595 PAD:9335 PAD:10179 0.026094
rPAD/1596 PAD:9335 PAD:10349 0.0222282
rPAD/1597 PAD:9335 PAD:15034 0.346154
rPAD/1598 PAD:9334 PAD:9336 0.0241118
rPAD/1599 PAD:9334 PAD:9335 0.346154
rPAD/1600 PAD:9332 PAD:9334 0.00419336
rPAD/1601 PAD:9331 PAD:9332 0.0241118
rPAD/1602 PAD:9330 PAD:10009 0.0294765
rPAD/1603 PAD:9330 PAD:10179 0.0188456
rPAD/1604 PAD:9330 PAD:15030 0.346154
rPAD/1605 PAD:9329 PAD:9331 0.0204426
rPAD/1606 PAD:9329 PAD:9330 0.346154
rPAD/1607 PAD:9327 PAD:9329 0.0319744
rPAD/1608 PAD:9326 PAD:9839 0.0328591
rPAD/1609 PAD:9326 PAD:10009 0.0154631
rPAD/1610 PAD:9326 PAD:15026 0.346154
rPAD/1611 PAD:9325 PAD:9327 0.0167734
rPAD/1612 PAD:9325 PAD:9326 0.346154
rPAD/1613 PAD:9323 PAD:9325 0.0356436
rPAD/1614 PAD:9321 PAD:9323 0.0293535
rPAD/1615 PAD:9321 PAD:15021 0.346154
rPAD/1616 PAD:9319 PAD:9321 0.0230635
rPAD/1617 PAD:9317 PAD:9319 0.0256843
rPAD/1618 PAD:9317 PAD:15017 0.346154
rPAD/1619 PAD:9314 PAD:9317 0.0487478
rPAD/1620 PAD:9314 PAD:15014 0.346154
rPAD/1621 PAD:9304 PAD:15000 0.0243668
rPAD/1622 PAD:9304 PAD:15004 0.9
rPAD/1623 PAD:9300 PAD:14598 0.0239738
rPAD/1624 PAD:9299 PAD:9300 1.5
rPAD/1625 PAD:9297 PAD:14992 0.0638646
rPAD/1626 PAD:9297 PAD:9300 0.0243668
rPAD/1627 PAD:9296 PAD:9299 0.0279
rPAD/1628 PAD:9296 PAD:9297 1.5
rPAD/1629 PAD:9293 PAD:9296 0.073125
rPAD/1630 PAD:9293 PAD:14992 1.5
rPAD/1631 PAD:9291 PAD:14989 0.00962882
rPAD/1632 PAD:9291 PAD:14992 0.0279039
rPAD/1633 PAD:9290 PAD:9293 0.03195
rPAD/1634 PAD:9290 PAD:9291 1.5
rPAD/1635 PAD:9288 PAD:9290 0.011025
rPAD/1636 PAD:9287 PAD:14987 0.0279039
rPAD/1637 PAD:9286 PAD:9288 0.052875
rPAD/1638 PAD:9286 PAD:9287 1.5
rPAD/1639 PAD:9284 PAD:14983 0.00451965
rPAD/1640 PAD:9284 PAD:9287 0.0279039
rPAD/1641 PAD:9283 PAD:9286 0.03195
rPAD/1642 PAD:9283 PAD:9284 1.5
rPAD/1643 PAD:9281 PAD:9283 0.005175
rPAD/1644 PAD:9280 PAD:14978 0.0273144
rPAD/1645 PAD:9280 PAD:14981 0.0279039
rPAD/1646 PAD:9279 PAD:9281 0.058725
rPAD/1647 PAD:9279 PAD:9280 1.5
rPAD/1648 PAD:9277 PAD:9279 0.031275
rPAD/1649 PAD:9276 PAD:14978 0.00058952
rPAD/1650 PAD:9275 PAD:9277 0.000675
rPAD/1651 PAD:9275 PAD:9276 1.5
rPAD/1652 PAD:9273 PAD:14973 0.0222052
rPAD/1653 PAD:9273 PAD:9276 0.0558079
rPAD/1654 PAD:9272 PAD:9275 0.0639
rPAD/1655 PAD:9272 PAD:9273 1.5
rPAD/1656 PAD:9270 PAD:9272 0.025425
rPAD/1657 PAD:9268 PAD:9270 0.006525
rPAD/1658 PAD:9268 PAD:14971 1.5
rPAD/1659 PAD:9265 PAD:9268 0.0639
rPAD/1660 PAD:9265 PAD:14968 1.5
rPAD/1661 PAD:9263 PAD:9265 0.019575
rPAD/1662 PAD:9262 PAD:14963 0.0558079
rPAD/1663 PAD:9262 PAD:14966 0.0108079
rPAD/1664 PAD:9261 PAD:9263 0.012375
rPAD/1665 PAD:9261 PAD:9262 1.5
rPAD/1666 PAD:9258 PAD:9261 0.0639
rPAD/1667 PAD:9258 PAD:14963 1.5
rPAD/1668 PAD:9256 PAD:9258 0.013725
rPAD/1669 PAD:9255 PAD:14958 0.0279039
rPAD/1670 PAD:9255 PAD:14961 0.015917
rPAD/1671 PAD:9254 PAD:9256 0.018225
rPAD/1672 PAD:9254 PAD:9255 1.5
rPAD/1673 PAD:9252 PAD:14955 0.00687773
rPAD/1674 PAD:9252 PAD:14958 0.0279039
rPAD/1675 PAD:9251 PAD:9254 0.0639
rPAD/1676 PAD:9251 PAD:9252 1.5
rPAD/1677 PAD:9249 PAD:9251 0.007875
rPAD/1678 PAD:9248 PAD:14952 0.0279039
rPAD/1679 PAD:9248 PAD:14955 0.0210262
rPAD/1680 PAD:9247 PAD:9249 0.024075
rPAD/1681 PAD:9247 PAD:9248 1.5
rPAD/1682 PAD:9245 PAD:14949 0.00176856
rPAD/1683 PAD:9245 PAD:14952 0.0279039
rPAD/1684 PAD:9244 PAD:9247 0.0639
rPAD/1685 PAD:9244 PAD:9245 1.5
rPAD/1686 PAD:9242 PAD:9244 0.002025
rPAD/1687 PAD:9240 PAD:9242 0.029925
rPAD/1688 PAD:9240 PAD:14947 1.5
rPAD/1689 PAD:9238 PAD:9240 0.060075
rPAD/1690 PAD:9237 PAD:14942 0.0279039
rPAD/1691 PAD:9237 PAD:14945 0.00334061
rPAD/1692 PAD:9236 PAD:9238 0.003825
rPAD/1693 PAD:9236 PAD:9237 1.5
rPAD/1694 PAD:9233 PAD:9236 0.03195
rPAD/1695 PAD:9233 PAD:14942 1.5
rPAD/1696 PAD:9231 PAD:9233 0.054225
rPAD/1697 PAD:9229 PAD:9231 0.009675
rPAD/1698 PAD:9229 PAD:14938 1.5
rPAD/1699 PAD:9227 PAD:14935 0.0422489
rPAD/1700 PAD:9227 PAD:14938 0.0279039
rPAD/1701 PAD:9226 PAD:9229 0.03195
rPAD/1702 PAD:9226 PAD:9227 1.5
rPAD/1703 PAD:9224 PAD:9226 0.048375
rPAD/1704 PAD:9222 PAD:9224 0.015525
rPAD/1705 PAD:9222 PAD:14933 1.5
rPAD/1706 PAD:9220 PAD:14929 0.0279039
rPAD/1707 PAD:9220 PAD:14933 0.0279039
rPAD/1708 PAD:9219 PAD:9222 0.03195
rPAD/1709 PAD:9219 PAD:9220 1.5
rPAD/1710 PAD:9217 PAD:9219 0.042525
rPAD/1711 PAD:9216 PAD:14927 0.0186681
rPAD/1712 PAD:9215 PAD:9217 0.021375
rPAD/1713 PAD:9215 PAD:9216 1.5
rPAD/1714 PAD:9213 PAD:14923 0.0279039
rPAD/1715 PAD:9213 PAD:9216 0.0279039
rPAD/1716 PAD:9212 PAD:9215 0.03195
rPAD/1717 PAD:9212 PAD:9213 1.5
rPAD/1718 PAD:9210 PAD:9212 0.036675
rPAD/1719 PAD:9209 PAD:14921 0.0237773
rPAD/1720 PAD:9208 PAD:9210 0.027225
rPAD/1721 PAD:9208 PAD:9209 1.5
rPAD/1722 PAD:9206 PAD:14916 0.0269214
rPAD/1723 PAD:9206 PAD:9209 0.0279039
rPAD/1724 PAD:9205 PAD:9208 0.03195
rPAD/1725 PAD:9205 PAD:9206 1.5
rPAD/1726 PAD:9203 PAD:9205 0.030825
rPAD/1727 PAD:9202 PAD:14913 0.0279039
rPAD/1728 PAD:9202 PAD:14916 0.0288865
rPAD/1729 PAD:9201 PAD:9203 0.033075
rPAD/1730 PAD:9201 PAD:9202 1.5
rPAD/1731 PAD:9198 PAD:9201 0.03195
rPAD/1732 PAD:9198 PAD:14913 1.5
rPAD/1733 PAD:9196 PAD:9198 0.024975
rPAD/1734 PAD:9194 PAD:9196 0.038925
rPAD/1735 PAD:9194 PAD:14909 1.5
rPAD/1736 PAD:9192 PAD:14906 0.0167031
rPAD/1737 PAD:9192 PAD:14909 0.0279039
rPAD/1738 PAD:9191 PAD:9194 0.03195
rPAD/1739 PAD:9191 PAD:9192 1.5
rPAD/1740 PAD:9189 PAD:9191 0.019125
rPAD/1741 PAD:9187 PAD:9189 0.044775
rPAD/1742 PAD:9187 PAD:14904 1.5
rPAD/1743 PAD:9185 PAD:14901 0.0115939
rPAD/1744 PAD:9185 PAD:14904 0.0279039
rPAD/1745 PAD:9184 PAD:9187 0.03195
rPAD/1746 PAD:9184 PAD:9185 1.5
rPAD/1747 PAD:9182 PAD:9184 0.013275
rPAD/1748 PAD:9181 PAD:14899 0.0279039
rPAD/1749 PAD:9180 PAD:9182 0.050625
rPAD/1750 PAD:9180 PAD:9181 1.5
rPAD/1751 PAD:9178 PAD:14895 0.00648472
rPAD/1752 PAD:9178 PAD:9181 0.0279039
rPAD/1753 PAD:9177 PAD:9180 0.03195
rPAD/1754 PAD:9177 PAD:9178 1.5
rPAD/1755 PAD:9175 PAD:9177 0.007425
rPAD/1756 PAD:9174 PAD:14889 0.0279039
rPAD/1757 PAD:9174 PAD:14893 0.0279039
rPAD/1758 PAD:9173 PAD:9175 0.056475
rPAD/1759 PAD:9173 PAD:9174 1.5
rPAD/1760 PAD:9170 PAD:9173 0.03195
rPAD/1761 PAD:9170 PAD:14889 1.5
rPAD/1762 PAD:9168 PAD:9170 0.001575
rPAD/1763 PAD:9167 PAD:14885 0.0241703
rPAD/1764 PAD:9167 PAD:14887 0.0544323
rPAD/1765 PAD:9166 PAD:9168 0.062325
rPAD/1766 PAD:9166 PAD:9167 1.5
rPAD/1767 PAD:9164 PAD:9166 0.027675
rPAD/1768 PAD:9162 PAD:9164 0.004275
rPAD/1769 PAD:9162 PAD:14883 1.5
rPAD/1770 PAD:9159 PAD:9162 0.0639
rPAD/1771 PAD:9159 PAD:14880 1.5
rPAD/1772 PAD:9157 PAD:9159 0.021825
rPAD/1773 PAD:9156 PAD:14875 0.0558079
rPAD/1774 PAD:9156 PAD:14878 0.0088428
rPAD/1775 PAD:9155 PAD:9157 0.010125
rPAD/1776 PAD:9155 PAD:9156 1.5
rPAD/1777 PAD:9152 PAD:9155 0.0639
rPAD/1778 PAD:9152 PAD:14875 1.5
rPAD/1779 PAD:9150 PAD:9152 0.015975
rPAD/1780 PAD:9149 PAD:14870 0.0279039
rPAD/1781 PAD:9149 PAD:14873 0.013952
rPAD/1782 PAD:9148 PAD:9150 0.015975
rPAD/1783 PAD:9148 PAD:9149 1.5
rPAD/1784 PAD:9146 PAD:14867 0.0088428
rPAD/1785 PAD:9146 PAD:14870 0.0279039
rPAD/1786 PAD:9145 PAD:9148 0.0639
rPAD/1787 PAD:9145 PAD:9146 1.5
rPAD/1788 PAD:9143 PAD:9145 0.010125
rPAD/1789 PAD:9142 PAD:14864 0.0279039
rPAD/1790 PAD:9142 PAD:14867 0.0190611
rPAD/1791 PAD:9141 PAD:9143 0.021825
rPAD/1792 PAD:9141 PAD:9142 1.5
rPAD/1793 PAD:9139 PAD:14861 0.00373362
rPAD/1794 PAD:9139 PAD:14864 0.0279039
rPAD/1795 PAD:9138 PAD:9141 0.0639
rPAD/1796 PAD:9138 PAD:9139 1.5
rPAD/1797 PAD:9136 PAD:9138 0.004275
rPAD/1798 PAD:9135 PAD:14857 0.0544323
rPAD/1799 PAD:9135 PAD:14861 0.0241703
rPAD/1800 PAD:9135 PAD:14860 0.9
rPAD/1801 PAD:9134 PAD:9136 0.027675
rPAD/1802 PAD:9134 PAD:9135 1.5
rPAD/1803 PAD:9132 PAD:9134 0.062325
rPAD/1804 PAD:9131 PAD:14857 0.00137555
rPAD/1805 PAD:9130 PAD:9132 0.001575
rPAD/1806 PAD:9130 PAD:9131 1.5
rPAD/1807 PAD:9128 PAD:14852 0.0493231
rPAD/1808 PAD:9128 PAD:9131 0.0279039
rPAD/1809 PAD:9128 PAD:14855 0.9
rPAD/1810 PAD:9127 PAD:9130 0.03195
rPAD/1811 PAD:9127 PAD:9128 1.5
rPAD/1812 PAD:9125 PAD:9127 0.056475
rPAD/1813 PAD:9123 PAD:9125 0.007425
rPAD/1814 PAD:9123 PAD:14850 1.5
rPAD/1815 PAD:9121 PAD:14847 0.044214
rPAD/1816 PAD:9121 PAD:14850 0.0279039
rPAD/1817 PAD:9120 PAD:9123 0.03195
rPAD/1818 PAD:9120 PAD:9121 1.5
rPAD/1819 PAD:9118 PAD:9120 0.050625
rPAD/1820 PAD:9116 PAD:9118 0.013275
rPAD/1821 PAD:9116 PAD:14845 1.5
rPAD/1822 PAD:9114 PAD:14841 0.0279039
rPAD/1823 PAD:9114 PAD:14845 0.0279039
rPAD/1824 PAD:9113 PAD:9116 0.03195
rPAD/1825 PAD:9113 PAD:9114 1.5
rPAD/1826 PAD:9111 PAD:9113 0.044775
rPAD/1827 PAD:9110 PAD:14839 0.0167031
rPAD/1828 PAD:9109 PAD:9111 0.019125
rPAD/1829 PAD:9109 PAD:9110 1.5
rPAD/1830 PAD:9107 PAD:14835 0.0279039
rPAD/1831 PAD:9107 PAD:9110 0.0279039
rPAD/1832 PAD:9106 PAD:9109 0.03195
rPAD/1833 PAD:9106 PAD:9107 1.5
rPAD/1834 PAD:9104 PAD:9106 0.038925
rPAD/1835 PAD:9103 PAD:14833 0.0218122
rPAD/1836 PAD:9102 PAD:9104 0.024975
rPAD/1837 PAD:9102 PAD:9103 1.5
rPAD/1838 PAD:9100 PAD:9103 0.0279039
rPAD/1839 PAD:9100 PAD:14831 0.9
rPAD/1840 PAD:9099 PAD:9102 0.03195
rPAD/1841 PAD:9099 PAD:9100 1.5
rPAD/1842 PAD:9097 PAD:9100 0.0279039
rPAD/1843 PAD:9096 PAD:9099 0.03195
rPAD/1844 PAD:9096 PAD:9097 1.5
rPAD/1845 PAD:9094 PAD:9450 0.0224017
rPAD/1846 PAD:9094 PAD:9097 0.0646507
rPAD/1847 PAD:9094 PAD:14827 0.9
rPAD/1848 PAD:9093 PAD:9096 0.074025
rPAD/1849 PAD:9093 PAD:9094 1.5
rPAD/1850 PAD:9090 PAD:14822 0.0243668
rPAD/1851 PAD:9089 PAD:9090 1.5
rPAD/1852 PAD:9086 PAD:9090 0.0243668
rPAD/1853 PAD:9086 PAD:9089 1.5279
rPAD/1854 PAD:9083 PAD:14599 0.0152215
rPAD/1855 PAD:9083 PAD:9449 0.0140134
rPAD/1856 PAD:9082 PAD:9083 2.25
rPAD/1857 PAD:9080 PAD:14599 0.012825
rPAD/1858 PAD:9079 PAD:9082 0.01395
rPAD/1859 PAD:9079 PAD:9080 0.586956
rPAD/1860 PAD:9077 PAD:9080 0.01395
rPAD/1861 PAD:9077 PAD:14814 0.225
rPAD/1862 PAD:9076 PAD:9079 0.01395
rPAD/1863 PAD:9076 PAD:9077 0.586956
rPAD/1864 PAD:9074 PAD:9077 0.0279
rPAD/1865 PAD:9074 PAD:14811 0.586956
rPAD/1866 PAD:9073 PAD:9076 0.0279
rPAD/1867 PAD:9073 PAD:9074 0.586956
rPAD/1868 PAD:9071 PAD:14806 0.01395
rPAD/1869 PAD:9071 PAD:9074 0.01395
rPAD/1870 PAD:9070 PAD:9073 0.01395
rPAD/1871 PAD:9070 PAD:9071 0.586956
rPAD/1872 PAD:9067 PAD:9070 0.0279
rPAD/1873 PAD:9067 PAD:14803 0.586956
rPAD/1874 PAD:9065 PAD:14799 0.01395
rPAD/1875 PAD:9065 PAD:14803 0.01395
rPAD/1876 PAD:9064 PAD:9067 0.01395
rPAD/1877 PAD:9064 PAD:9065 0.586956
rPAD/1878 PAD:9062 PAD:14795 0.01395
rPAD/1879 PAD:9062 PAD:14799 0.01395
rPAD/1880 PAD:9061 PAD:9064 0.0279
rPAD/1881 PAD:9061 PAD:9062 0.586956
rPAD/1882 PAD:9058 PAD:9061 0.0279
rPAD/1883 PAD:9058 PAD:14792 0.586956
rPAD/1884 PAD:9056 PAD:14788 0.01395
rPAD/1885 PAD:9056 PAD:14792 0.01395
rPAD/1886 PAD:9055 PAD:9058 0.01395
rPAD/1887 PAD:9055 PAD:9056 0.586956
rPAD/1888 PAD:9052 PAD:9055 0.0279
rPAD/1889 PAD:9052 PAD:14785 0.586956
rPAD/1890 PAD:9049 PAD:9052 0.01395
rPAD/1891 PAD:9049 PAD:14782 0.586956
rPAD/1892 PAD:9047 PAD:14778 0.01395
rPAD/1893 PAD:9047 PAD:14782 0.01395
rPAD/1894 PAD:9046 PAD:9049 0.01395
rPAD/1895 PAD:9046 PAD:9047 0.586956
rPAD/1896 PAD:9044 PAD:14774 0.01395
rPAD/1897 PAD:9044 PAD:14778 0.01395
rPAD/1898 PAD:9043 PAD:9046 0.0279
rPAD/1899 PAD:9043 PAD:9044 0.586956
rPAD/1900 PAD:9040 PAD:9043 0.0279
rPAD/1901 PAD:9040 PAD:14771 0.586956
rPAD/1902 PAD:9038 PAD:14767 0.01395
rPAD/1903 PAD:9038 PAD:14771 0.01395
rPAD/1904 PAD:9037 PAD:9040 0.01395
rPAD/1905 PAD:9037 PAD:9038 0.586956
rPAD/1906 PAD:9034 PAD:9037 0.0279
rPAD/1907 PAD:9034 PAD:14764 0.586956
rPAD/1908 PAD:9032 PAD:14760 0.01395
rPAD/1909 PAD:9032 PAD:14764 0.01395
rPAD/1910 PAD:9031 PAD:9034 0.01395
rPAD/1911 PAD:9031 PAD:9032 0.586956
rPAD/1912 PAD:9029 PAD:14760 0.01395
rPAD/1913 PAD:9029 PAD:14758 0.586956
rPAD/1914 PAD:9028 PAD:9031 0.0279
rPAD/1915 PAD:9028 PAD:9029 0.586956
rPAD/1916 PAD:9026 PAD:14753 0.01395
rPAD/1917 PAD:9026 PAD:9029 0.01395
rPAD/1918 PAD:9025 PAD:9028 0.01395
rPAD/1919 PAD:9025 PAD:9026 0.586956
rPAD/1920 PAD:9022 PAD:9025 0.0279
rPAD/1921 PAD:9022 PAD:14750 0.586956
rPAD/1922 PAD:9020 PAD:14746 0.01395
rPAD/1923 PAD:9020 PAD:14750 0.01395
rPAD/1924 PAD:9019 PAD:9022 0.01395
rPAD/1925 PAD:9019 PAD:9020 0.586956
rPAD/1926 PAD:9017 PAD:14742 0.01395
rPAD/1927 PAD:9017 PAD:14746 0.01395
rPAD/1928 PAD:9016 PAD:9019 0.0279
rPAD/1929 PAD:9016 PAD:9017 0.586956
rPAD/1930 PAD:9013 PAD:9016 0.0279
rPAD/1931 PAD:9013 PAD:14739 0.586956
rPAD/1932 PAD:9011 PAD:14735 0.01395
rPAD/1933 PAD:9011 PAD:14739 0.01395
rPAD/1934 PAD:9010 PAD:9013 0.01395
rPAD/1935 PAD:9010 PAD:9011 0.586956
rPAD/1936 PAD:9007 PAD:9010 0.0279
rPAD/1937 PAD:9007 PAD:14732 0.586956
rPAD/1938 PAD:9004 PAD:9007 0.01395
rPAD/1939 PAD:9004 PAD:14729 0.586956
rPAD/1940 PAD:9002 PAD:14725 0.01395
rPAD/1941 PAD:9002 PAD:14729 0.01395
rPAD/1942 PAD:9001 PAD:9004 0.01395
rPAD/1943 PAD:9001 PAD:9002 0.586956
rPAD/1944 PAD:8999 PAD:14721 0.01395
rPAD/1945 PAD:8999 PAD:14725 0.01395
rPAD/1946 PAD:8998 PAD:9001 0.0279
rPAD/1947 PAD:8998 PAD:8999 0.586956
rPAD/1948 PAD:8995 PAD:8998 0.0279
rPAD/1949 PAD:8995 PAD:14718 0.586956
rPAD/1950 PAD:8993 PAD:14714 0.01395
rPAD/1951 PAD:8993 PAD:14718 0.01395
rPAD/1952 PAD:8992 PAD:8995 0.01395
rPAD/1953 PAD:8992 PAD:8993 0.586956
rPAD/1954 PAD:8989 PAD:8992 0.0279
rPAD/1955 PAD:8989 PAD:14711 0.586956
rPAD/1956 PAD:8987 PAD:14707 0.01395
rPAD/1957 PAD:8987 PAD:14711 0.01395
rPAD/1958 PAD:8986 PAD:8989 0.01395
rPAD/1959 PAD:8986 PAD:8987 0.586956
rPAD/1960 PAD:8984 PAD:14707 0.01395
rPAD/1961 PAD:8983 PAD:8986 0.0279
rPAD/1962 PAD:8983 PAD:8984 0.586956
rPAD/1963 PAD:8981 PAD:14700 0.01395
rPAD/1964 PAD:8981 PAD:8984 0.01395
rPAD/1965 PAD:8980 PAD:8983 0.01395
rPAD/1966 PAD:8980 PAD:8981 0.586956
rPAD/1967 PAD:8977 PAD:8980 0.0279
rPAD/1968 PAD:8977 PAD:14697 0.586956
rPAD/1969 PAD:8975 PAD:14693 0.01395
rPAD/1970 PAD:8975 PAD:14697 0.01395
rPAD/1971 PAD:8974 PAD:8977 0.01395
rPAD/1972 PAD:8974 PAD:8975 0.586956
rPAD/1973 PAD:8972 PAD:14689 0.01395
rPAD/1974 PAD:8972 PAD:14693 0.01395
rPAD/1975 PAD:8971 PAD:8974 0.0279
rPAD/1976 PAD:8971 PAD:8972 0.586956
rPAD/1977 PAD:8968 PAD:8971 0.0279
rPAD/1978 PAD:8968 PAD:14686 0.586956
rPAD/1979 PAD:8966 PAD:14682 0.01395
rPAD/1980 PAD:8966 PAD:14686 0.01395
rPAD/1981 PAD:8965 PAD:8968 0.01395
rPAD/1982 PAD:8965 PAD:8966 0.586956
rPAD/1983 PAD:8962 PAD:8965 0.0279
rPAD/1984 PAD:8962 PAD:14679 0.586956
rPAD/1985 PAD:8959 PAD:8962 0.01395
rPAD/1986 PAD:8959 PAD:14676 0.586956
rPAD/1987 PAD:8957 PAD:14672 0.01395
rPAD/1988 PAD:8957 PAD:14676 0.01395
rPAD/1989 PAD:8956 PAD:8959 0.01395
rPAD/1990 PAD:8956 PAD:8957 0.586956
rPAD/1991 PAD:8954 PAD:14668 0.01395
rPAD/1992 PAD:8954 PAD:14672 0.01395
rPAD/1993 PAD:8953 PAD:8956 0.0279
rPAD/1994 PAD:8953 PAD:8954 0.586956
rPAD/1995 PAD:8950 PAD:8953 0.0279
rPAD/1996 PAD:8950 PAD:14665 0.586956
rPAD/1997 PAD:8948 PAD:14661 0.01395
rPAD/1998 PAD:8948 PAD:14665 0.01395
rPAD/1999 PAD:8947 PAD:8950 0.01395
rPAD/2000 PAD:8947 PAD:8948 0.586956
rPAD/2001 PAD:8944 PAD:8947 0.0279
rPAD/2002 PAD:8944 PAD:14658 0.586956
rPAD/2003 PAD:8942 PAD:14654 0.01395
rPAD/2004 PAD:8942 PAD:14658 0.01395
rPAD/2005 PAD:8941 PAD:8944 0.01395
rPAD/2006 PAD:8941 PAD:8942 0.586956
rPAD/2007 PAD:8939 PAD:14654 0.01395
rPAD/2008 PAD:8938 PAD:8941 0.0279
rPAD/2009 PAD:8938 PAD:8939 0.586956
rPAD/2010 PAD:8936 PAD:14647 0.01395
rPAD/2011 PAD:8936 PAD:8939 0.01395
rPAD/2012 PAD:8935 PAD:8938 0.01395
rPAD/2013 PAD:8935 PAD:8936 0.586956
rPAD/2014 PAD:8932 PAD:8935 0.0279
rPAD/2015 PAD:8932 PAD:14644 0.586956
rPAD/2016 PAD:8930 PAD:14640 0.01395
rPAD/2017 PAD:8930 PAD:14644 0.01395
rPAD/2018 PAD:8929 PAD:8932 0.01395
rPAD/2019 PAD:8929 PAD:8930 0.586956
rPAD/2020 PAD:8927 PAD:14636 0.01395
rPAD/2021 PAD:8927 PAD:14640 0.01395
rPAD/2022 PAD:8926 PAD:8929 0.0279
rPAD/2023 PAD:8926 PAD:8927 0.586956
rPAD/2024 PAD:8923 PAD:8926 0.0279
rPAD/2025 PAD:8923 PAD:14633 0.586956
rPAD/2026 PAD:8921 PAD:14629 0.01395
rPAD/2027 PAD:8921 PAD:14633 0.01395
rPAD/2028 PAD:8920 PAD:8923 0.01395
rPAD/2029 PAD:8920 PAD:8921 0.586956
rPAD/2030 PAD:8917 PAD:8920 0.0279
rPAD/2031 PAD:8917 PAD:14626 0.586956
rPAD/2032 PAD:8914 PAD:8917 0.01395
rPAD/2033 PAD:8914 PAD:14623 0.586956
rPAD/2034 PAD:8912 PAD:14619 0.01395
rPAD/2035 PAD:8912 PAD:14623 0.01395
rPAD/2036 PAD:8911 PAD:8914 0.01395
rPAD/2037 PAD:8911 PAD:8912 0.586956
rPAD/2038 PAD:8909 PAD:14615 0.01395
rPAD/2039 PAD:8909 PAD:14619 0.01395
rPAD/2040 PAD:8908 PAD:8911 0.0279
rPAD/2041 PAD:8908 PAD:8909 0.586956
rPAD/2042 PAD:8905 PAD:8908 0.0279
rPAD/2043 PAD:8905 PAD:14612 0.586956
rPAD/2044 PAD:8903 PAD:14608 0.01395
rPAD/2045 PAD:8903 PAD:14612 0.01395
rPAD/2046 PAD:8902 PAD:8905 0.01395
rPAD/2047 PAD:8902 PAD:8903 0.586956
rPAD/2048 PAD:8899 PAD:8902 0.0279
rPAD/2049 PAD:8899 PAD:14605 0.586956
rPAD/2050 PAD:8897 PAD:14601 0.01395
rPAD/2051 PAD:8897 PAD:14605 0.01395
rPAD/2052 PAD:8896 PAD:8899 0.01395
rPAD/2053 PAD:8896 PAD:8897 0.586956
rPAD/2054 PAD:8893 PAD:8896 0.0279
rPAD/2055 PAD:8893 PAD:9297 0.586956
rPAD/2056 PAD:8891 PAD:9444 0.000786255
rPAD/2057 PAD:8891 PAD:9082 0.007875
rPAD/2058 PAD:8891 PAD:9449 1.53171
rPAD/2059 PAD:8890 PAD:9299 0.02745
rPAD/2060 PAD:8890 PAD:9304 1.15659
rPAD/2061 PAD:8890 PAD:8893 0.002925
rPAD/2062 PAD:8889 PAD:14429 0.0100588
rPAD/2063 PAD:8889 PAD:14597 1.5
rPAD/2064 PAD:8888 PAD:9439 0.0670908
rPAD/2065 PAD:8888 PAD:8889 1.5
rPAD/2066 PAD:8886 PAD:8889 0.0751765
rPAD/2067 PAD:8886 PAD:14594 1.5
rPAD/2068 PAD:8885 PAD:8888 0.0751765
rPAD/2069 PAD:8885 PAD:8886 1.5
rPAD/2070 PAD:8883 PAD:14587 0.0751765
rPAD/2071 PAD:8883 PAD:8886 0.0375882
rPAD/2072 PAD:8883 PAD:14591 1.5
rPAD/2073 PAD:8882 PAD:8885 0.0375882
rPAD/2074 PAD:8882 PAD:8883 1.5
rPAD/2075 PAD:8879 PAD:8882 0.0751765
rPAD/2076 PAD:8879 PAD:14587 1.5
rPAD/2077 PAD:8877 PAD:14587 0.0375882
rPAD/2078 PAD:8877 PAD:14585 1.5
rPAD/2079 PAD:8876 PAD:8879 0.0375882
rPAD/2080 PAD:8876 PAD:8877 1.5
rPAD/2081 PAD:8874 PAD:8877 0.0751765
rPAD/2082 PAD:8874 PAD:14582 1.5
rPAD/2083 PAD:8873 PAD:8876 0.0751765
rPAD/2084 PAD:8873 PAD:8874 1.5
rPAD/2085 PAD:8871 PAD:8874 0.0375882
rPAD/2086 PAD:8871 PAD:14579 1.5
rPAD/2087 PAD:8870 PAD:8873 0.0375882
rPAD/2088 PAD:8870 PAD:8871 1.5
rPAD/2089 PAD:8868 PAD:8871 0.0751765
rPAD/2090 PAD:8868 PAD:14576 1.5
rPAD/2091 PAD:8867 PAD:8870 0.0751765
rPAD/2092 PAD:8867 PAD:8868 1.5
rPAD/2093 PAD:8865 PAD:8868 0.0375882
rPAD/2094 PAD:8865 PAD:14573 1.5
rPAD/2095 PAD:8864 PAD:8867 0.0375882
rPAD/2096 PAD:8864 PAD:8865 1.5
rPAD/2097 PAD:8862 PAD:8865 0.0751765
rPAD/2098 PAD:8862 PAD:14570 1.5
rPAD/2099 PAD:8861 PAD:8864 0.0751765
rPAD/2100 PAD:8861 PAD:8862 1.5
rPAD/2101 PAD:8859 PAD:8862 0.0375882
rPAD/2102 PAD:8859 PAD:14567 1.5
rPAD/2103 PAD:8858 PAD:8861 0.0375882
rPAD/2104 PAD:8858 PAD:8859 1.5
rPAD/2105 PAD:8856 PAD:8859 0.0751765
rPAD/2106 PAD:8856 PAD:14564 1.5
rPAD/2107 PAD:8855 PAD:8858 0.0751765
rPAD/2108 PAD:8855 PAD:8856 1.5
rPAD/2109 PAD:8853 PAD:8856 0.0375882
rPAD/2110 PAD:8853 PAD:14561 1.5
rPAD/2111 PAD:8852 PAD:8855 0.0375882
rPAD/2112 PAD:8852 PAD:8853 1.5
rPAD/2113 PAD:8850 PAD:8853 0.0751765
rPAD/2114 PAD:8850 PAD:14558 1.5
rPAD/2115 PAD:8849 PAD:8852 0.0751765
rPAD/2116 PAD:8849 PAD:8850 1.5
rPAD/2117 PAD:8847 PAD:14551 0.0751765
rPAD/2118 PAD:8847 PAD:8850 0.0375882
rPAD/2119 PAD:8847 PAD:14555 1.5
rPAD/2120 PAD:8846 PAD:8849 0.0375882
rPAD/2121 PAD:8846 PAD:8847 1.5
rPAD/2122 PAD:8843 PAD:8846 0.0751765
rPAD/2123 PAD:8843 PAD:14551 1.5
rPAD/2124 PAD:8841 PAD:14545 0.0751765
rPAD/2125 PAD:8841 PAD:14551 0.0375882
rPAD/2126 PAD:8841 PAD:14549 1.5
rPAD/2127 PAD:8840 PAD:8843 0.0375882
rPAD/2128 PAD:8840 PAD:8841 1.5
rPAD/2129 PAD:8837 PAD:8840 0.0751765
rPAD/2130 PAD:8837 PAD:14545 1.5
rPAD/2131 PAD:8834 PAD:8837 0.0375882
rPAD/2132 PAD:8834 PAD:14542 1.5
rPAD/2133 PAD:8831 PAD:8834 0.0751765
rPAD/2134 PAD:8831 PAD:14539 1.5
rPAD/2135 PAD:8829 PAD:14533 0.0751765
rPAD/2136 PAD:8829 PAD:14539 0.0375882
rPAD/2137 PAD:8829 PAD:14537 1.5
rPAD/2138 PAD:8828 PAD:8831 0.0375882
rPAD/2139 PAD:8828 PAD:8829 1.5
rPAD/2140 PAD:8825 PAD:8828 0.0751765
rPAD/2141 PAD:8825 PAD:14533 1.5
rPAD/2142 PAD:8822 PAD:8825 0.0375882
rPAD/2143 PAD:8822 PAD:14530 1.5
rPAD/2144 PAD:8820 PAD:14530 0.0751765
rPAD/2145 PAD:8820 PAD:14528 1.5
rPAD/2146 PAD:8819 PAD:8822 0.0751765
rPAD/2147 PAD:8819 PAD:8820 1.5
rPAD/2148 PAD:8817 PAD:8820 0.0375882
rPAD/2149 PAD:8817 PAD:14525 1.5
rPAD/2150 PAD:8816 PAD:8819 0.0375882
rPAD/2151 PAD:8816 PAD:8817 1.5
rPAD/2152 PAD:8814 PAD:8817 0.0751765
rPAD/2153 PAD:8814 PAD:14522 1.5
rPAD/2154 PAD:8813 PAD:8816 0.0751765
rPAD/2155 PAD:8813 PAD:8814 1.5
rPAD/2156 PAD:8811 PAD:8814 0.0375882
rPAD/2157 PAD:8811 PAD:14519 1.5
rPAD/2158 PAD:8810 PAD:8813 0.0375882
rPAD/2159 PAD:8810 PAD:8811 1.5
rPAD/2160 PAD:8808 PAD:8811 0.0751765
rPAD/2161 PAD:8808 PAD:14516 1.5
rPAD/2162 PAD:8807 PAD:8810 0.0751765
rPAD/2163 PAD:8807 PAD:8808 1.5
rPAD/2164 PAD:8805 PAD:14509 0.0751765
rPAD/2165 PAD:8805 PAD:8808 0.0375882
rPAD/2166 PAD:8805 PAD:14513 1.5
rPAD/2167 PAD:8804 PAD:8807 0.0375882
rPAD/2168 PAD:8804 PAD:8805 1.5
rPAD/2169 PAD:8801 PAD:8804 0.0751765
rPAD/2170 PAD:8801 PAD:14509 1.5
rPAD/2171 PAD:8799 PAD:14509 0.0375882
rPAD/2172 PAD:8799 PAD:14507 1.5
rPAD/2173 PAD:8798 PAD:8801 0.0375882
rPAD/2174 PAD:8798 PAD:8799 1.5
rPAD/2175 PAD:8796 PAD:8799 0.0751765
rPAD/2176 PAD:8796 PAD:14504 1.5
rPAD/2177 PAD:8795 PAD:8798 0.0751765
rPAD/2178 PAD:8795 PAD:8796 1.5
rPAD/2179 PAD:8793 PAD:14497 0.0751765
rPAD/2180 PAD:8793 PAD:8796 0.0375882
rPAD/2181 PAD:8793 PAD:14501 1.5
rPAD/2182 PAD:8792 PAD:8795 0.0375882
rPAD/2183 PAD:8792 PAD:8793 1.5
rPAD/2184 PAD:8789 PAD:8792 0.0751765
rPAD/2185 PAD:8789 PAD:14497 1.5
rPAD/2186 PAD:8786 PAD:8789 0.0375882
rPAD/2187 PAD:8786 PAD:14494 1.5
rPAD/2188 PAD:8783 PAD:8786 0.0751765
rPAD/2189 PAD:8783 PAD:14491 1.5
rPAD/2190 PAD:8780 PAD:8783 0.0375882
rPAD/2191 PAD:8780 PAD:14488 1.5
rPAD/2192 PAD:8777 PAD:8780 0.0751765
rPAD/2193 PAD:8777 PAD:14485 1.5
rPAD/2194 PAD:8775 PAD:14485 0.0375882
rPAD/2195 PAD:8775 PAD:14483 1.5
rPAD/2196 PAD:8774 PAD:8777 0.0375882
rPAD/2197 PAD:8774 PAD:8775 1.5
rPAD/2198 PAD:8772 PAD:14476 0.0375882
rPAD/2199 PAD:8772 PAD:8775 0.0751765
rPAD/2200 PAD:8772 PAD:14480 1.5
rPAD/2201 PAD:8771 PAD:8774 0.0751765
rPAD/2202 PAD:8771 PAD:8772 1.5
rPAD/2203 PAD:8768 PAD:8771 0.0375882
rPAD/2204 PAD:8768 PAD:14476 1.5
rPAD/2205 PAD:8766 PAD:14476 0.0751765
rPAD/2206 PAD:8766 PAD:14474 1.5
rPAD/2207 PAD:8765 PAD:8768 0.0751765
rPAD/2208 PAD:8765 PAD:8766 1.5
rPAD/2209 PAD:8763 PAD:8766 0.0375882
rPAD/2210 PAD:8763 PAD:14471 1.5
rPAD/2211 PAD:8762 PAD:8765 0.0375882
rPAD/2212 PAD:8762 PAD:8763 1.5
rPAD/2213 PAD:8760 PAD:8763 0.0751765
rPAD/2214 PAD:8760 PAD:14468 1.5
rPAD/2215 PAD:8759 PAD:8762 0.0751765
rPAD/2216 PAD:8759 PAD:8760 1.5
rPAD/2217 PAD:8757 PAD:8760 0.0375882
rPAD/2218 PAD:8757 PAD:14465 1.5
rPAD/2219 PAD:8756 PAD:8759 0.0375882
rPAD/2220 PAD:8756 PAD:8757 1.5
rPAD/2221 PAD:8754 PAD:8757 0.0751765
rPAD/2222 PAD:8754 PAD:14462 1.5
rPAD/2223 PAD:8753 PAD:8756 0.0751765
rPAD/2224 PAD:8753 PAD:8754 1.5
rPAD/2225 PAD:8751 PAD:14455 0.0751765
rPAD/2226 PAD:8751 PAD:8754 0.0375882
rPAD/2227 PAD:8751 PAD:14459 1.5
rPAD/2228 PAD:8750 PAD:8753 0.0375882
rPAD/2229 PAD:8750 PAD:8751 1.5
rPAD/2230 PAD:8747 PAD:8750 0.0751765
rPAD/2231 PAD:8747 PAD:14455 1.5
rPAD/2232 PAD:8745 PAD:14455 0.0375882
rPAD/2233 PAD:8745 PAD:14453 1.5
rPAD/2234 PAD:8744 PAD:8747 0.0375882
rPAD/2235 PAD:8744 PAD:8745 1.5
rPAD/2236 PAD:8742 PAD:8745 0.0751765
rPAD/2237 PAD:8742 PAD:14450 1.5
rPAD/2238 PAD:8741 PAD:8744 0.0751765
rPAD/2239 PAD:8741 PAD:8742 1.5
rPAD/2240 PAD:8739 PAD:8742 0.0375882
rPAD/2241 PAD:8739 PAD:14447 1.5
rPAD/2242 PAD:8738 PAD:8741 0.0375882
rPAD/2243 PAD:8738 PAD:8739 1.5
rPAD/2244 PAD:8736 PAD:8739 0.0751765
rPAD/2245 PAD:8736 PAD:14444 1.5
rPAD/2246 PAD:8735 PAD:8738 0.0751765
rPAD/2247 PAD:8735 PAD:8736 1.5
rPAD/2248 PAD:8733 PAD:8736 0.0375882
rPAD/2249 PAD:8733 PAD:14441 1.5
rPAD/2250 PAD:8732 PAD:8735 0.0375882
rPAD/2251 PAD:8732 PAD:8733 1.5
rPAD/2252 PAD:8730 PAD:8733 0.0751765
rPAD/2253 PAD:8730 PAD:14438 1.5
rPAD/2254 PAD:8729 PAD:8732 0.0751765
rPAD/2255 PAD:8729 PAD:8730 1.5
rPAD/2256 PAD:8727 PAD:8730 0.0375882
rPAD/2257 PAD:8727 PAD:14435 1.5
rPAD/2258 PAD:8726 PAD:8729 0.0375882
rPAD/2259 PAD:8726 PAD:8727 1.5
rPAD/2260 PAD:8724 PAD:14989 0.0283817
rPAD/2261 PAD:8724 PAD:8727 0.0751765
rPAD/2262 PAD:8724 PAD:14432 1.5
rPAD/2263 PAD:8723 PAD:9288 0.0378785
rPAD/2264 PAD:8723 PAD:8726 0.0751765
rPAD/2265 PAD:8723 PAD:8724 1.5
rPAD/2266 PAD:8719 PAD:14259 0.0100588
rPAD/2267 PAD:8719 PAD:14427 1.5
rPAD/2268 PAD:8718 PAD:9435 0.0670908
rPAD/2269 PAD:8718 PAD:8719 1.5
rPAD/2270 PAD:8716 PAD:8719 0.0751765
rPAD/2271 PAD:8716 PAD:14424 1.5
rPAD/2272 PAD:8715 PAD:8718 0.0751765
rPAD/2273 PAD:8715 PAD:8716 1.5
rPAD/2274 PAD:8713 PAD:14417 0.0751765
rPAD/2275 PAD:8713 PAD:8716 0.0375882
rPAD/2276 PAD:8713 PAD:14421 1.5
rPAD/2277 PAD:8712 PAD:8715 0.0375882
rPAD/2278 PAD:8712 PAD:8713 1.5
rPAD/2279 PAD:8709 PAD:8712 0.0751765
rPAD/2280 PAD:8709 PAD:14417 1.5
rPAD/2281 PAD:8707 PAD:14417 0.0375882
rPAD/2282 PAD:8707 PAD:14415 1.5
rPAD/2283 PAD:8706 PAD:8709 0.0375882
rPAD/2284 PAD:8706 PAD:8707 1.5
rPAD/2285 PAD:8704 PAD:8707 0.0751765
rPAD/2286 PAD:8704 PAD:14412 1.5
rPAD/2287 PAD:8703 PAD:8706 0.0751765
rPAD/2288 PAD:8703 PAD:8704 1.5
rPAD/2289 PAD:8701 PAD:8704 0.0375882
rPAD/2290 PAD:8701 PAD:14409 1.5
rPAD/2291 PAD:8700 PAD:8703 0.0375882
rPAD/2292 PAD:8700 PAD:8701 1.5
rPAD/2293 PAD:8698 PAD:8701 0.0751765
rPAD/2294 PAD:8698 PAD:14406 1.5
rPAD/2295 PAD:8697 PAD:8700 0.0751765
rPAD/2296 PAD:8697 PAD:8698 1.5
rPAD/2297 PAD:8695 PAD:8698 0.0375882
rPAD/2298 PAD:8695 PAD:14403 1.5
rPAD/2299 PAD:8694 PAD:8697 0.0375882
rPAD/2300 PAD:8694 PAD:8695 1.5
rPAD/2301 PAD:8692 PAD:8695 0.0751765
rPAD/2302 PAD:8692 PAD:14400 1.5
rPAD/2303 PAD:8691 PAD:8694 0.0751765
rPAD/2304 PAD:8691 PAD:8692 1.5
rPAD/2305 PAD:8689 PAD:8692 0.0375882
rPAD/2306 PAD:8689 PAD:14397 1.5
rPAD/2307 PAD:8688 PAD:8691 0.0375882
rPAD/2308 PAD:8688 PAD:8689 1.5
rPAD/2309 PAD:8686 PAD:8689 0.0751765
rPAD/2310 PAD:8686 PAD:14394 1.5
rPAD/2311 PAD:8685 PAD:8688 0.0751765
rPAD/2312 PAD:8685 PAD:8686 1.5
rPAD/2313 PAD:8683 PAD:8686 0.0375882
rPAD/2314 PAD:8683 PAD:14391 1.5
rPAD/2315 PAD:8682 PAD:8685 0.0375882
rPAD/2316 PAD:8682 PAD:8683 1.5
rPAD/2317 PAD:8680 PAD:8683 0.0751765
rPAD/2318 PAD:8680 PAD:14388 1.5
rPAD/2319 PAD:8679 PAD:8682 0.0751765
rPAD/2320 PAD:8679 PAD:8680 1.5
rPAD/2321 PAD:8677 PAD:14381 0.0751765
rPAD/2322 PAD:8677 PAD:8680 0.0375882
rPAD/2323 PAD:8677 PAD:14385 1.5
rPAD/2324 PAD:8676 PAD:8679 0.0375882
rPAD/2325 PAD:8676 PAD:8677 1.5
rPAD/2326 PAD:8673 PAD:8676 0.0751765
rPAD/2327 PAD:8673 PAD:14381 1.5
rPAD/2328 PAD:8671 PAD:14375 0.0751765
rPAD/2329 PAD:8671 PAD:14381 0.0375882
rPAD/2330 PAD:8671 PAD:14379 1.5
rPAD/2331 PAD:8670 PAD:8673 0.0375882
rPAD/2332 PAD:8670 PAD:8671 1.5
rPAD/2333 PAD:8667 PAD:8670 0.0751765
rPAD/2334 PAD:8667 PAD:14375 1.5
rPAD/2335 PAD:8664 PAD:8667 0.0375882
rPAD/2336 PAD:8664 PAD:14372 1.5
rPAD/2337 PAD:8661 PAD:8664 0.0751765
rPAD/2338 PAD:8661 PAD:14369 1.5
rPAD/2339 PAD:8659 PAD:14363 0.0751765
rPAD/2340 PAD:8659 PAD:14369 0.0375882
rPAD/2341 PAD:8659 PAD:14367 1.5
rPAD/2342 PAD:8658 PAD:8661 0.0375882
rPAD/2343 PAD:8658 PAD:8659 1.5
rPAD/2344 PAD:8655 PAD:8658 0.0751765
rPAD/2345 PAD:8655 PAD:14363 1.5
rPAD/2346 PAD:8652 PAD:8655 0.0375882
rPAD/2347 PAD:8652 PAD:14360 1.5
rPAD/2348 PAD:8650 PAD:14360 0.0751765
rPAD/2349 PAD:8650 PAD:14358 1.5
rPAD/2350 PAD:8649 PAD:8652 0.0751765
rPAD/2351 PAD:8649 PAD:8650 1.5
rPAD/2352 PAD:8647 PAD:8650 0.0375882
rPAD/2353 PAD:8647 PAD:14355 1.5
rPAD/2354 PAD:8646 PAD:8649 0.0375882
rPAD/2355 PAD:8646 PAD:8647 1.5
rPAD/2356 PAD:8644 PAD:8647 0.0751765
rPAD/2357 PAD:8644 PAD:14352 1.5
rPAD/2358 PAD:8643 PAD:8646 0.0751765
rPAD/2359 PAD:8643 PAD:8644 1.5
rPAD/2360 PAD:8641 PAD:8644 0.0375882
rPAD/2361 PAD:8641 PAD:14349 1.5
rPAD/2362 PAD:8640 PAD:8643 0.0375882
rPAD/2363 PAD:8640 PAD:8641 1.5
rPAD/2364 PAD:8638 PAD:8641 0.0751765
rPAD/2365 PAD:8638 PAD:14346 1.5
rPAD/2366 PAD:8637 PAD:8640 0.0751765
rPAD/2367 PAD:8637 PAD:8638 1.5
rPAD/2368 PAD:8635 PAD:14339 0.0751765
rPAD/2369 PAD:8635 PAD:8638 0.0375882
rPAD/2370 PAD:8635 PAD:14343 1.5
rPAD/2371 PAD:8634 PAD:8637 0.0375882
rPAD/2372 PAD:8634 PAD:8635 1.5
rPAD/2373 PAD:8631 PAD:8634 0.0751765
rPAD/2374 PAD:8631 PAD:14339 1.5
rPAD/2375 PAD:8629 PAD:14339 0.0375882
rPAD/2376 PAD:8629 PAD:14337 1.5
rPAD/2377 PAD:8628 PAD:8631 0.0375882
rPAD/2378 PAD:8628 PAD:8629 1.5
rPAD/2379 PAD:8626 PAD:8629 0.0751765
rPAD/2380 PAD:8626 PAD:14334 1.5
rPAD/2381 PAD:8625 PAD:8628 0.0751765
rPAD/2382 PAD:8625 PAD:8626 1.5
rPAD/2383 PAD:8623 PAD:14327 0.0751765
rPAD/2384 PAD:8623 PAD:8626 0.0375882
rPAD/2385 PAD:8623 PAD:14331 1.5
rPAD/2386 PAD:8622 PAD:8625 0.0375882
rPAD/2387 PAD:8622 PAD:8623 1.5
rPAD/2388 PAD:8619 PAD:8622 0.0751765
rPAD/2389 PAD:8619 PAD:14327 1.5
rPAD/2390 PAD:8616 PAD:8619 0.0375882
rPAD/2391 PAD:8616 PAD:14324 1.5
rPAD/2392 PAD:8613 PAD:8616 0.0751765
rPAD/2393 PAD:8613 PAD:14321 1.5
rPAD/2394 PAD:8610 PAD:8613 0.0375882
rPAD/2395 PAD:8610 PAD:14318 1.5
rPAD/2396 PAD:8607 PAD:8610 0.0751765
rPAD/2397 PAD:8607 PAD:14315 1.5
rPAD/2398 PAD:8605 PAD:14315 0.0375882
rPAD/2399 PAD:8605 PAD:14313 1.5
rPAD/2400 PAD:8604 PAD:8607 0.0375882
rPAD/2401 PAD:8604 PAD:8605 1.5
rPAD/2402 PAD:8602 PAD:14306 0.0375882
rPAD/2403 PAD:8602 PAD:8605 0.0751765
rPAD/2404 PAD:8602 PAD:14310 1.5
rPAD/2405 PAD:8601 PAD:8604 0.0751765
rPAD/2406 PAD:8601 PAD:8602 1.5
rPAD/2407 PAD:8598 PAD:8601 0.0375882
rPAD/2408 PAD:8598 PAD:14306 1.5
rPAD/2409 PAD:8596 PAD:14306 0.0751765
rPAD/2410 PAD:8596 PAD:14304 1.5
rPAD/2411 PAD:8595 PAD:8598 0.0751765
rPAD/2412 PAD:8595 PAD:8596 1.5
rPAD/2413 PAD:8593 PAD:8596 0.0375882
rPAD/2414 PAD:8593 PAD:14301 1.5
rPAD/2415 PAD:8592 PAD:8595 0.0375882
rPAD/2416 PAD:8592 PAD:8593 1.5
rPAD/2417 PAD:8590 PAD:8593 0.0751765
rPAD/2418 PAD:8590 PAD:14298 1.5
rPAD/2419 PAD:8589 PAD:8592 0.0751765
rPAD/2420 PAD:8589 PAD:8590 1.5
rPAD/2421 PAD:8587 PAD:8590 0.0375882
rPAD/2422 PAD:8587 PAD:14295 1.5
rPAD/2423 PAD:8586 PAD:8589 0.0375882
rPAD/2424 PAD:8586 PAD:8587 1.5
rPAD/2425 PAD:8584 PAD:8587 0.0751765
rPAD/2426 PAD:8584 PAD:14292 1.5
rPAD/2427 PAD:8583 PAD:8586 0.0751765
rPAD/2428 PAD:8583 PAD:8584 1.5
rPAD/2429 PAD:8581 PAD:14285 0.0751765
rPAD/2430 PAD:8581 PAD:8584 0.0375882
rPAD/2431 PAD:8581 PAD:14289 1.5
rPAD/2432 PAD:8580 PAD:8583 0.0375882
rPAD/2433 PAD:8580 PAD:8581 1.5
rPAD/2434 PAD:8577 PAD:8580 0.0751765
rPAD/2435 PAD:8577 PAD:14285 1.5
rPAD/2436 PAD:8575 PAD:14285 0.0375882
rPAD/2437 PAD:8575 PAD:14283 1.5
rPAD/2438 PAD:8574 PAD:8577 0.0375882
rPAD/2439 PAD:8574 PAD:8575 1.5
rPAD/2440 PAD:8572 PAD:8575 0.0751765
rPAD/2441 PAD:8572 PAD:14280 1.5
rPAD/2442 PAD:8571 PAD:8574 0.0751765
rPAD/2443 PAD:8571 PAD:8572 1.5
rPAD/2444 PAD:8569 PAD:8572 0.0375882
rPAD/2445 PAD:8569 PAD:14277 1.5
rPAD/2446 PAD:8568 PAD:8571 0.0375882
rPAD/2447 PAD:8568 PAD:8569 1.5
rPAD/2448 PAD:8566 PAD:8569 0.0751765
rPAD/2449 PAD:8566 PAD:14274 1.5
rPAD/2450 PAD:8565 PAD:8568 0.0751765
rPAD/2451 PAD:8565 PAD:8566 1.5
rPAD/2452 PAD:8563 PAD:8566 0.0375882
rPAD/2453 PAD:8563 PAD:14271 1.5
rPAD/2454 PAD:8562 PAD:8565 0.0375882
rPAD/2455 PAD:8562 PAD:8563 1.5
rPAD/2456 PAD:8560 PAD:8563 0.0751765
rPAD/2457 PAD:8560 PAD:14268 1.5
rPAD/2458 PAD:8559 PAD:8562 0.0751765
rPAD/2459 PAD:8559 PAD:8560 1.5
rPAD/2460 PAD:8557 PAD:8560 0.0375882
rPAD/2461 PAD:8557 PAD:14265 1.5
rPAD/2462 PAD:8556 PAD:8559 0.0375882
rPAD/2463 PAD:8556 PAD:8557 1.5
rPAD/2464 PAD:8554 PAD:14983 0.0283817
rPAD/2465 PAD:8554 PAD:8557 0.0751765
rPAD/2466 PAD:8554 PAD:14262 1.5
rPAD/2467 PAD:8553 PAD:9281 0.0378785
rPAD/2468 PAD:8553 PAD:8556 0.0751765
rPAD/2469 PAD:8553 PAD:8554 1.5
rPAD/2470 PAD:8549 PAD:14089 0.0100588
rPAD/2471 PAD:8549 PAD:14257 1.5
rPAD/2472 PAD:8548 PAD:9431 0.0670908
rPAD/2473 PAD:8548 PAD:8549 1.5
rPAD/2474 PAD:8546 PAD:8549 0.0751765
rPAD/2475 PAD:8546 PAD:14254 1.5
rPAD/2476 PAD:8545 PAD:8548 0.0751765
rPAD/2477 PAD:8545 PAD:8546 1.5
rPAD/2478 PAD:8543 PAD:14247 0.0751765
rPAD/2479 PAD:8543 PAD:8546 0.0375882
rPAD/2480 PAD:8543 PAD:14251 1.5
rPAD/2481 PAD:8542 PAD:8545 0.0375882
rPAD/2482 PAD:8542 PAD:8543 1.5
rPAD/2483 PAD:8539 PAD:8542 0.0751765
rPAD/2484 PAD:8539 PAD:14247 1.5
rPAD/2485 PAD:8537 PAD:14247 0.0375882
rPAD/2486 PAD:8537 PAD:14245 1.5
rPAD/2487 PAD:8536 PAD:8539 0.0375882
rPAD/2488 PAD:8536 PAD:8537 1.5
rPAD/2489 PAD:8534 PAD:8537 0.0751765
rPAD/2490 PAD:8534 PAD:14242 1.5
rPAD/2491 PAD:8533 PAD:8536 0.0751765
rPAD/2492 PAD:8533 PAD:8534 1.5
rPAD/2493 PAD:8531 PAD:8534 0.0375882
rPAD/2494 PAD:8531 PAD:14239 1.5
rPAD/2495 PAD:8530 PAD:8533 0.0375882
rPAD/2496 PAD:8530 PAD:8531 1.5
rPAD/2497 PAD:8528 PAD:8531 0.0751765
rPAD/2498 PAD:8528 PAD:14236 1.5
rPAD/2499 PAD:8527 PAD:8530 0.0751765
rPAD/2500 PAD:8527 PAD:8528 1.5
rPAD/2501 PAD:8525 PAD:8528 0.0375882
rPAD/2502 PAD:8525 PAD:14233 1.5
rPAD/2503 PAD:8524 PAD:8527 0.0375882
rPAD/2504 PAD:8524 PAD:8525 1.5
rPAD/2505 PAD:8522 PAD:8525 0.0751765
rPAD/2506 PAD:8522 PAD:14230 1.5
rPAD/2507 PAD:8521 PAD:8524 0.0751765
rPAD/2508 PAD:8521 PAD:8522 1.5
rPAD/2509 PAD:8519 PAD:8522 0.0375882
rPAD/2510 PAD:8519 PAD:14227 1.5
rPAD/2511 PAD:8518 PAD:8521 0.0375882
rPAD/2512 PAD:8518 PAD:8519 1.5
rPAD/2513 PAD:8516 PAD:8519 0.0751765
rPAD/2514 PAD:8516 PAD:14224 1.5
rPAD/2515 PAD:8515 PAD:8518 0.0751765
rPAD/2516 PAD:8515 PAD:8516 1.5
rPAD/2517 PAD:8513 PAD:8516 0.0375882
rPAD/2518 PAD:8513 PAD:14221 1.5
rPAD/2519 PAD:8512 PAD:8515 0.0375882
rPAD/2520 PAD:8512 PAD:8513 1.5
rPAD/2521 PAD:8510 PAD:8513 0.0751765
rPAD/2522 PAD:8510 PAD:14218 1.5
rPAD/2523 PAD:8509 PAD:8512 0.0751765
rPAD/2524 PAD:8509 PAD:8510 1.5
rPAD/2525 PAD:8507 PAD:14211 0.0751765
rPAD/2526 PAD:8507 PAD:8510 0.0375882
rPAD/2527 PAD:8507 PAD:14215 1.5
rPAD/2528 PAD:8506 PAD:8509 0.0375882
rPAD/2529 PAD:8506 PAD:8507 1.5
rPAD/2530 PAD:8503 PAD:8506 0.0751765
rPAD/2531 PAD:8503 PAD:14211 1.5
rPAD/2532 PAD:8501 PAD:14205 0.0751765
rPAD/2533 PAD:8501 PAD:14211 0.0375882
rPAD/2534 PAD:8501 PAD:14209 1.5
rPAD/2535 PAD:8500 PAD:8503 0.0375882
rPAD/2536 PAD:8500 PAD:8501 1.5
rPAD/2537 PAD:8497 PAD:8500 0.0751765
rPAD/2538 PAD:8497 PAD:14205 1.5
rPAD/2539 PAD:8494 PAD:8497 0.0375882
rPAD/2540 PAD:8494 PAD:14202 1.5
rPAD/2541 PAD:8491 PAD:8494 0.0751765
rPAD/2542 PAD:8491 PAD:14199 1.5
rPAD/2543 PAD:8489 PAD:14193 0.0751765
rPAD/2544 PAD:8489 PAD:14199 0.0375882
rPAD/2545 PAD:8489 PAD:14197 1.5
rPAD/2546 PAD:8488 PAD:8491 0.0375882
rPAD/2547 PAD:8488 PAD:8489 1.5
rPAD/2548 PAD:8485 PAD:8488 0.0751765
rPAD/2549 PAD:8485 PAD:14193 1.5
rPAD/2550 PAD:8482 PAD:8485 0.0375882
rPAD/2551 PAD:8482 PAD:14190 1.5
rPAD/2552 PAD:8480 PAD:14190 0.0751765
rPAD/2553 PAD:8480 PAD:14188 1.5
rPAD/2554 PAD:8479 PAD:8482 0.0751765
rPAD/2555 PAD:8479 PAD:8480 1.5
rPAD/2556 PAD:8477 PAD:8480 0.0375882
rPAD/2557 PAD:8477 PAD:14185 1.5
rPAD/2558 PAD:8476 PAD:8479 0.0375882
rPAD/2559 PAD:8476 PAD:8477 1.5
rPAD/2560 PAD:8474 PAD:8477 0.0751765
rPAD/2561 PAD:8474 PAD:14182 1.5
rPAD/2562 PAD:8473 PAD:8476 0.0751765
rPAD/2563 PAD:8473 PAD:8474 1.5
rPAD/2564 PAD:8471 PAD:8474 0.0375882
rPAD/2565 PAD:8471 PAD:14179 1.5
rPAD/2566 PAD:8470 PAD:8473 0.0375882
rPAD/2567 PAD:8470 PAD:8471 1.5
rPAD/2568 PAD:8468 PAD:8471 0.0751765
rPAD/2569 PAD:8468 PAD:14176 1.5
rPAD/2570 PAD:8467 PAD:8470 0.0751765
rPAD/2571 PAD:8467 PAD:8468 1.5
rPAD/2572 PAD:8465 PAD:14169 0.0751765
rPAD/2573 PAD:8465 PAD:8468 0.0375882
rPAD/2574 PAD:8465 PAD:14173 1.5
rPAD/2575 PAD:8464 PAD:8467 0.0375882
rPAD/2576 PAD:8464 PAD:8465 1.5
rPAD/2577 PAD:8461 PAD:8464 0.0751765
rPAD/2578 PAD:8461 PAD:14169 1.5
rPAD/2579 PAD:8459 PAD:14169 0.0375882
rPAD/2580 PAD:8459 PAD:14167 1.5
rPAD/2581 PAD:8458 PAD:8461 0.0375882
rPAD/2582 PAD:8458 PAD:8459 1.5
rPAD/2583 PAD:8456 PAD:8459 0.0751765
rPAD/2584 PAD:8456 PAD:14164 1.5
rPAD/2585 PAD:8455 PAD:8458 0.0751765
rPAD/2586 PAD:8455 PAD:8456 1.5
rPAD/2587 PAD:8453 PAD:14157 0.0751765
rPAD/2588 PAD:8453 PAD:8456 0.0375882
rPAD/2589 PAD:8453 PAD:14161 1.5
rPAD/2590 PAD:8452 PAD:8455 0.0375882
rPAD/2591 PAD:8452 PAD:8453 1.5
rPAD/2592 PAD:8449 PAD:8452 0.0751765
rPAD/2593 PAD:8449 PAD:14157 1.5
rPAD/2594 PAD:8446 PAD:8449 0.0375882
rPAD/2595 PAD:8446 PAD:14154 1.5
rPAD/2596 PAD:8443 PAD:8446 0.0751765
rPAD/2597 PAD:8443 PAD:14151 1.5
rPAD/2598 PAD:8440 PAD:8443 0.0375882
rPAD/2599 PAD:8440 PAD:14148 1.5
rPAD/2600 PAD:8437 PAD:8440 0.0751765
rPAD/2601 PAD:8437 PAD:14145 1.5
rPAD/2602 PAD:8435 PAD:14145 0.0375882
rPAD/2603 PAD:8435 PAD:14143 1.5
rPAD/2604 PAD:8434 PAD:8437 0.0375882
rPAD/2605 PAD:8434 PAD:8435 1.5
rPAD/2606 PAD:8432 PAD:14136 0.0375882
rPAD/2607 PAD:8432 PAD:8435 0.0751765
rPAD/2608 PAD:8432 PAD:14140 1.5
rPAD/2609 PAD:8431 PAD:8434 0.0751765
rPAD/2610 PAD:8431 PAD:8432 1.5
rPAD/2611 PAD:8428 PAD:8431 0.0375882
rPAD/2612 PAD:8428 PAD:14136 1.5
rPAD/2613 PAD:8426 PAD:14136 0.0751765
rPAD/2614 PAD:8426 PAD:14134 1.5
rPAD/2615 PAD:8425 PAD:8428 0.0751765
rPAD/2616 PAD:8425 PAD:8426 1.5
rPAD/2617 PAD:8423 PAD:8426 0.0375882
rPAD/2618 PAD:8423 PAD:14131 1.5
rPAD/2619 PAD:8422 PAD:8425 0.0375882
rPAD/2620 PAD:8422 PAD:8423 1.5
rPAD/2621 PAD:8420 PAD:8423 0.0751765
rPAD/2622 PAD:8420 PAD:14128 1.5
rPAD/2623 PAD:8419 PAD:8422 0.0751765
rPAD/2624 PAD:8419 PAD:8420 1.5
rPAD/2625 PAD:8417 PAD:8420 0.0375882
rPAD/2626 PAD:8417 PAD:14125 1.5
rPAD/2627 PAD:8416 PAD:8419 0.0375882
rPAD/2628 PAD:8416 PAD:8417 1.5
rPAD/2629 PAD:8414 PAD:8417 0.0751765
rPAD/2630 PAD:8414 PAD:14122 1.5
rPAD/2631 PAD:8413 PAD:8416 0.0751765
rPAD/2632 PAD:8413 PAD:8414 1.5
rPAD/2633 PAD:8411 PAD:14115 0.0751765
rPAD/2634 PAD:8411 PAD:8414 0.0375882
rPAD/2635 PAD:8411 PAD:14119 1.5
rPAD/2636 PAD:8410 PAD:8413 0.0375882
rPAD/2637 PAD:8410 PAD:8411 1.5
rPAD/2638 PAD:8407 PAD:8410 0.0751765
rPAD/2639 PAD:8407 PAD:14115 1.5
rPAD/2640 PAD:8405 PAD:14115 0.0375882
rPAD/2641 PAD:8405 PAD:14113 1.5
rPAD/2642 PAD:8404 PAD:8407 0.0375882
rPAD/2643 PAD:8404 PAD:8405 1.5
rPAD/2644 PAD:8402 PAD:8405 0.0751765
rPAD/2645 PAD:8402 PAD:14110 1.5
rPAD/2646 PAD:8401 PAD:8404 0.0751765
rPAD/2647 PAD:8401 PAD:8402 1.5
rPAD/2648 PAD:8399 PAD:8402 0.0375882
rPAD/2649 PAD:8399 PAD:14107 1.5
rPAD/2650 PAD:8398 PAD:8401 0.0375882
rPAD/2651 PAD:8398 PAD:8399 1.5
rPAD/2652 PAD:8396 PAD:8399 0.0751765
rPAD/2653 PAD:8396 PAD:14104 1.5
rPAD/2654 PAD:8395 PAD:8398 0.0751765
rPAD/2655 PAD:8395 PAD:8396 1.5
rPAD/2656 PAD:8393 PAD:8396 0.0375882
rPAD/2657 PAD:8393 PAD:14101 1.5
rPAD/2658 PAD:8392 PAD:8395 0.0375882
rPAD/2659 PAD:8392 PAD:8393 1.5
rPAD/2660 PAD:8390 PAD:8393 0.0751765
rPAD/2661 PAD:8390 PAD:14098 1.5
rPAD/2662 PAD:8389 PAD:8392 0.0751765
rPAD/2663 PAD:8389 PAD:8390 1.5
rPAD/2664 PAD:8387 PAD:8390 0.0375882
rPAD/2665 PAD:8387 PAD:14095 1.5
rPAD/2666 PAD:8386 PAD:8389 0.0375882
rPAD/2667 PAD:8386 PAD:8387 1.5
rPAD/2668 PAD:8384 PAD:14978 0.0283817
rPAD/2669 PAD:8384 PAD:8387 0.0751765
rPAD/2670 PAD:8384 PAD:14092 1.5
rPAD/2671 PAD:8383 PAD:9277 0.0378785
rPAD/2672 PAD:8383 PAD:8386 0.0751765
rPAD/2673 PAD:8383 PAD:8384 1.5
rPAD/2674 PAD:8379 PAD:13919 0.0100588
rPAD/2675 PAD:8379 PAD:14087 1.5
rPAD/2676 PAD:8378 PAD:9427 0.0670908
rPAD/2677 PAD:8378 PAD:8379 1.5
rPAD/2678 PAD:8376 PAD:8379 0.0751765
rPAD/2679 PAD:8376 PAD:14084 1.5
rPAD/2680 PAD:8375 PAD:8378 0.0751765
rPAD/2681 PAD:8375 PAD:8376 1.5
rPAD/2682 PAD:8373 PAD:14077 0.0751765
rPAD/2683 PAD:8373 PAD:8376 0.0375882
rPAD/2684 PAD:8373 PAD:14081 1.5
rPAD/2685 PAD:8372 PAD:8375 0.0375882
rPAD/2686 PAD:8372 PAD:8373 1.5
rPAD/2687 PAD:8369 PAD:8372 0.0751765
rPAD/2688 PAD:8369 PAD:14077 1.5
rPAD/2689 PAD:8367 PAD:14077 0.0375882
rPAD/2690 PAD:8367 PAD:14075 1.5
rPAD/2691 PAD:8366 PAD:8369 0.0375882
rPAD/2692 PAD:8366 PAD:8367 1.5
rPAD/2693 PAD:8364 PAD:8367 0.0751765
rPAD/2694 PAD:8364 PAD:14072 1.5
rPAD/2695 PAD:8363 PAD:8366 0.0751765
rPAD/2696 PAD:8363 PAD:8364 1.5
rPAD/2697 PAD:8361 PAD:8364 0.0375882
rPAD/2698 PAD:8361 PAD:14069 1.5
rPAD/2699 PAD:8360 PAD:8363 0.0375882
rPAD/2700 PAD:8360 PAD:8361 1.5
rPAD/2701 PAD:8358 PAD:8361 0.0751765
rPAD/2702 PAD:8358 PAD:14066 1.5
rPAD/2703 PAD:8357 PAD:8360 0.0751765
rPAD/2704 PAD:8357 PAD:8358 1.5
rPAD/2705 PAD:8355 PAD:8358 0.0375882
rPAD/2706 PAD:8355 PAD:14063 1.5
rPAD/2707 PAD:8354 PAD:8357 0.0375882
rPAD/2708 PAD:8354 PAD:8355 1.5
rPAD/2709 PAD:8352 PAD:8355 0.0751765
rPAD/2710 PAD:8352 PAD:14060 1.5
rPAD/2711 PAD:8351 PAD:8354 0.0751765
rPAD/2712 PAD:8351 PAD:8352 1.5
rPAD/2713 PAD:8349 PAD:8352 0.0375882
rPAD/2714 PAD:8349 PAD:14057 1.5
rPAD/2715 PAD:8348 PAD:8351 0.0375882
rPAD/2716 PAD:8348 PAD:8349 1.5
rPAD/2717 PAD:8346 PAD:8349 0.0751765
rPAD/2718 PAD:8346 PAD:14054 1.5
rPAD/2719 PAD:8345 PAD:8348 0.0751765
rPAD/2720 PAD:8345 PAD:8346 1.5
rPAD/2721 PAD:8343 PAD:8346 0.0375882
rPAD/2722 PAD:8343 PAD:14051 1.5
rPAD/2723 PAD:8342 PAD:8345 0.0375882
rPAD/2724 PAD:8342 PAD:8343 1.5
rPAD/2725 PAD:8340 PAD:8343 0.0751765
rPAD/2726 PAD:8340 PAD:14048 1.5
rPAD/2727 PAD:8339 PAD:8342 0.0751765
rPAD/2728 PAD:8339 PAD:8340 1.5
rPAD/2729 PAD:8337 PAD:14041 0.0751765
rPAD/2730 PAD:8337 PAD:8340 0.0375882
rPAD/2731 PAD:8337 PAD:14045 1.5
rPAD/2732 PAD:8336 PAD:8339 0.0375882
rPAD/2733 PAD:8336 PAD:8337 1.5
rPAD/2734 PAD:8333 PAD:8336 0.0751765
rPAD/2735 PAD:8333 PAD:14041 1.5
rPAD/2736 PAD:8331 PAD:14035 0.0751765
rPAD/2737 PAD:8331 PAD:14041 0.0375882
rPAD/2738 PAD:8331 PAD:14039 1.5
rPAD/2739 PAD:8330 PAD:8333 0.0375882
rPAD/2740 PAD:8330 PAD:8331 1.5
rPAD/2741 PAD:8327 PAD:8330 0.0751765
rPAD/2742 PAD:8327 PAD:14035 1.5
rPAD/2743 PAD:8324 PAD:8327 0.0375882
rPAD/2744 PAD:8324 PAD:14032 1.5
rPAD/2745 PAD:8321 PAD:8324 0.0751765
rPAD/2746 PAD:8321 PAD:14029 1.5
rPAD/2747 PAD:8319 PAD:14023 0.0751765
rPAD/2748 PAD:8319 PAD:14029 0.0375882
rPAD/2749 PAD:8319 PAD:14027 1.5
rPAD/2750 PAD:8318 PAD:8321 0.0375882
rPAD/2751 PAD:8318 PAD:8319 1.5
rPAD/2752 PAD:8315 PAD:8318 0.0751765
rPAD/2753 PAD:8315 PAD:14023 1.5
rPAD/2754 PAD:8312 PAD:8315 0.0375882
rPAD/2755 PAD:8312 PAD:14020 1.5
rPAD/2756 PAD:8310 PAD:14020 0.0751765
rPAD/2757 PAD:8310 PAD:14018 1.5
rPAD/2758 PAD:8309 PAD:8312 0.0751765
rPAD/2759 PAD:8309 PAD:8310 1.5
rPAD/2760 PAD:8307 PAD:8310 0.0375882
rPAD/2761 PAD:8307 PAD:14015 1.5
rPAD/2762 PAD:8306 PAD:8309 0.0375882
rPAD/2763 PAD:8306 PAD:8307 1.5
rPAD/2764 PAD:8304 PAD:8307 0.0751765
rPAD/2765 PAD:8304 PAD:14012 1.5
rPAD/2766 PAD:8303 PAD:8306 0.0751765
rPAD/2767 PAD:8303 PAD:8304 1.5
rPAD/2768 PAD:8301 PAD:8304 0.0375882
rPAD/2769 PAD:8301 PAD:14009 1.5
rPAD/2770 PAD:8300 PAD:8303 0.0375882
rPAD/2771 PAD:8300 PAD:8301 1.5
rPAD/2772 PAD:8298 PAD:8301 0.0751765
rPAD/2773 PAD:8298 PAD:14006 1.5
rPAD/2774 PAD:8297 PAD:8300 0.0751765
rPAD/2775 PAD:8297 PAD:8298 1.5
rPAD/2776 PAD:8295 PAD:13999 0.0751765
rPAD/2777 PAD:8295 PAD:8298 0.0375882
rPAD/2778 PAD:8295 PAD:14003 1.5
rPAD/2779 PAD:8294 PAD:8297 0.0375882
rPAD/2780 PAD:8294 PAD:8295 1.5
rPAD/2781 PAD:8291 PAD:8294 0.0751765
rPAD/2782 PAD:8291 PAD:13999 1.5
rPAD/2783 PAD:8289 PAD:13999 0.0375882
rPAD/2784 PAD:8289 PAD:13997 1.5
rPAD/2785 PAD:8288 PAD:8291 0.0375882
rPAD/2786 PAD:8288 PAD:8289 1.5
rPAD/2787 PAD:8286 PAD:8289 0.0751765
rPAD/2788 PAD:8286 PAD:13994 1.5
rPAD/2789 PAD:8285 PAD:8288 0.0751765
rPAD/2790 PAD:8285 PAD:8286 1.5
rPAD/2791 PAD:8283 PAD:13987 0.0751765
rPAD/2792 PAD:8283 PAD:8286 0.0375882
rPAD/2793 PAD:8283 PAD:13991 1.5
rPAD/2794 PAD:8282 PAD:8285 0.0375882
rPAD/2795 PAD:8282 PAD:8283 1.5
rPAD/2796 PAD:8279 PAD:8282 0.0751765
rPAD/2797 PAD:8279 PAD:13987 1.5
rPAD/2798 PAD:8276 PAD:8279 0.0375882
rPAD/2799 PAD:8276 PAD:13984 1.5
rPAD/2800 PAD:8273 PAD:8276 0.0751765
rPAD/2801 PAD:8273 PAD:13981 1.5
rPAD/2802 PAD:8270 PAD:8273 0.0375882
rPAD/2803 PAD:8270 PAD:13978 1.5
rPAD/2804 PAD:8267 PAD:8270 0.0751765
rPAD/2805 PAD:8267 PAD:13975 1.5
rPAD/2806 PAD:8265 PAD:13975 0.0375882
rPAD/2807 PAD:8265 PAD:13973 1.5
rPAD/2808 PAD:8264 PAD:8267 0.0375882
rPAD/2809 PAD:8264 PAD:8265 1.5
rPAD/2810 PAD:8262 PAD:13966 0.0375882
rPAD/2811 PAD:8262 PAD:8265 0.0751765
rPAD/2812 PAD:8262 PAD:13970 1.5
rPAD/2813 PAD:8261 PAD:8264 0.0751765
rPAD/2814 PAD:8261 PAD:8262 1.5
rPAD/2815 PAD:8258 PAD:8261 0.0375882
rPAD/2816 PAD:8258 PAD:13966 1.5
rPAD/2817 PAD:8256 PAD:13966 0.0751765
rPAD/2818 PAD:8256 PAD:13964 1.5
rPAD/2819 PAD:8255 PAD:8258 0.0751765
rPAD/2820 PAD:8255 PAD:8256 1.5
rPAD/2821 PAD:8253 PAD:8256 0.0375882
rPAD/2822 PAD:8253 PAD:13961 1.5
rPAD/2823 PAD:8252 PAD:8255 0.0375882
rPAD/2824 PAD:8252 PAD:8253 1.5
rPAD/2825 PAD:8250 PAD:8253 0.0751765
rPAD/2826 PAD:8250 PAD:13958 1.5
rPAD/2827 PAD:8249 PAD:8252 0.0751765
rPAD/2828 PAD:8249 PAD:8250 1.5
rPAD/2829 PAD:8247 PAD:8250 0.0375882
rPAD/2830 PAD:8247 PAD:13955 1.5
rPAD/2831 PAD:8246 PAD:8249 0.0375882
rPAD/2832 PAD:8246 PAD:8247 1.5
rPAD/2833 PAD:8244 PAD:8247 0.0751765
rPAD/2834 PAD:8244 PAD:13952 1.5
rPAD/2835 PAD:8243 PAD:8246 0.0751765
rPAD/2836 PAD:8243 PAD:8244 1.5
rPAD/2837 PAD:8241 PAD:13945 0.0751765
rPAD/2838 PAD:8241 PAD:8244 0.0375882
rPAD/2839 PAD:8241 PAD:13949 1.5
rPAD/2840 PAD:8240 PAD:8243 0.0375882
rPAD/2841 PAD:8240 PAD:8241 1.5
rPAD/2842 PAD:8237 PAD:8240 0.0751765
rPAD/2843 PAD:8237 PAD:13945 1.5
rPAD/2844 PAD:8235 PAD:13945 0.0375882
rPAD/2845 PAD:8235 PAD:13943 1.5
rPAD/2846 PAD:8234 PAD:8237 0.0375882
rPAD/2847 PAD:8234 PAD:8235 1.5
rPAD/2848 PAD:8232 PAD:8235 0.0751765
rPAD/2849 PAD:8232 PAD:13940 1.5
rPAD/2850 PAD:8231 PAD:8234 0.0751765
rPAD/2851 PAD:8231 PAD:8232 1.5
rPAD/2852 PAD:8229 PAD:8232 0.0375882
rPAD/2853 PAD:8229 PAD:13937 1.5
rPAD/2854 PAD:8228 PAD:8231 0.0375882
rPAD/2855 PAD:8228 PAD:8229 1.5
rPAD/2856 PAD:8226 PAD:8229 0.0751765
rPAD/2857 PAD:8226 PAD:13934 1.5
rPAD/2858 PAD:8225 PAD:8228 0.0751765
rPAD/2859 PAD:8225 PAD:8226 1.5
rPAD/2860 PAD:8223 PAD:8226 0.0375882
rPAD/2861 PAD:8223 PAD:13931 1.5
rPAD/2862 PAD:8222 PAD:8225 0.0375882
rPAD/2863 PAD:8222 PAD:8223 1.5
rPAD/2864 PAD:8220 PAD:8223 0.0751765
rPAD/2865 PAD:8220 PAD:13928 1.5
rPAD/2866 PAD:8219 PAD:8222 0.0751765
rPAD/2867 PAD:8219 PAD:8220 1.5
rPAD/2868 PAD:8217 PAD:8220 0.0375882
rPAD/2869 PAD:8217 PAD:13925 1.5
rPAD/2870 PAD:8216 PAD:8219 0.0375882
rPAD/2871 PAD:8216 PAD:8217 1.5
rPAD/2872 PAD:8214 PAD:14973 0.0283817
rPAD/2873 PAD:8214 PAD:8217 0.0751765
rPAD/2874 PAD:8214 PAD:13922 1.5
rPAD/2875 PAD:8213 PAD:9270 0.0378785
rPAD/2876 PAD:8213 PAD:8216 0.0751765
rPAD/2877 PAD:8213 PAD:8214 1.5
rPAD/2878 PAD:8209 PAD:13749 0.0100588
rPAD/2879 PAD:8209 PAD:13917 1.5
rPAD/2880 PAD:8208 PAD:9422 0.0670908
rPAD/2881 PAD:8208 PAD:8209 1.5
rPAD/2882 PAD:8206 PAD:8209 0.0751765
rPAD/2883 PAD:8206 PAD:13914 1.5
rPAD/2884 PAD:8205 PAD:8208 0.0751765
rPAD/2885 PAD:8205 PAD:8206 1.5
rPAD/2886 PAD:8203 PAD:13907 0.0751765
rPAD/2887 PAD:8203 PAD:8206 0.0375882
rPAD/2888 PAD:8203 PAD:13911 1.5
rPAD/2889 PAD:8202 PAD:8205 0.0375882
rPAD/2890 PAD:8202 PAD:8203 1.5
rPAD/2891 PAD:8199 PAD:8202 0.0751765
rPAD/2892 PAD:8199 PAD:13907 1.5
rPAD/2893 PAD:8197 PAD:13907 0.0375882
rPAD/2894 PAD:8197 PAD:13905 1.5
rPAD/2895 PAD:8196 PAD:8199 0.0375882
rPAD/2896 PAD:8196 PAD:8197 1.5
rPAD/2897 PAD:8194 PAD:8197 0.0751765
rPAD/2898 PAD:8194 PAD:13902 1.5
rPAD/2899 PAD:8193 PAD:8196 0.0751765
rPAD/2900 PAD:8193 PAD:8194 1.5
rPAD/2901 PAD:8191 PAD:8194 0.0375882
rPAD/2902 PAD:8191 PAD:13899 1.5
rPAD/2903 PAD:8190 PAD:8193 0.0375882
rPAD/2904 PAD:8190 PAD:8191 1.5
rPAD/2905 PAD:8188 PAD:8191 0.0751765
rPAD/2906 PAD:8188 PAD:13896 1.5
rPAD/2907 PAD:8187 PAD:8190 0.0751765
rPAD/2908 PAD:8187 PAD:8188 1.5
rPAD/2909 PAD:8185 PAD:8188 0.0375882
rPAD/2910 PAD:8185 PAD:13893 1.5
rPAD/2911 PAD:8184 PAD:8187 0.0375882
rPAD/2912 PAD:8184 PAD:8185 1.5
rPAD/2913 PAD:8182 PAD:8185 0.0751765
rPAD/2914 PAD:8182 PAD:13890 1.5
rPAD/2915 PAD:8181 PAD:8184 0.0751765
rPAD/2916 PAD:8181 PAD:8182 1.5
rPAD/2917 PAD:8179 PAD:8182 0.0375882
rPAD/2918 PAD:8179 PAD:13887 1.5
rPAD/2919 PAD:8178 PAD:8181 0.0375882
rPAD/2920 PAD:8178 PAD:8179 1.5
rPAD/2921 PAD:8176 PAD:8179 0.0751765
rPAD/2922 PAD:8176 PAD:13884 1.5
rPAD/2923 PAD:8175 PAD:8178 0.0751765
rPAD/2924 PAD:8175 PAD:8176 1.5
rPAD/2925 PAD:8173 PAD:8176 0.0375882
rPAD/2926 PAD:8173 PAD:13881 1.5
rPAD/2927 PAD:8172 PAD:8175 0.0375882
rPAD/2928 PAD:8172 PAD:8173 1.5
rPAD/2929 PAD:8170 PAD:8173 0.0751765
rPAD/2930 PAD:8170 PAD:13878 1.5
rPAD/2931 PAD:8169 PAD:8172 0.0751765
rPAD/2932 PAD:8169 PAD:8170 1.5
rPAD/2933 PAD:8167 PAD:13871 0.0751765
rPAD/2934 PAD:8167 PAD:8170 0.0375882
rPAD/2935 PAD:8167 PAD:13875 1.5
rPAD/2936 PAD:8166 PAD:8169 0.0375882
rPAD/2937 PAD:8166 PAD:8167 1.5
rPAD/2938 PAD:8163 PAD:8166 0.0751765
rPAD/2939 PAD:8163 PAD:13871 1.5
rPAD/2940 PAD:8161 PAD:13865 0.0751765
rPAD/2941 PAD:8161 PAD:13871 0.0375882
rPAD/2942 PAD:8161 PAD:13869 1.5
rPAD/2943 PAD:8160 PAD:8163 0.0375882
rPAD/2944 PAD:8160 PAD:8161 1.5
rPAD/2945 PAD:8157 PAD:8160 0.0751765
rPAD/2946 PAD:8157 PAD:13865 1.5
rPAD/2947 PAD:8154 PAD:8157 0.0375882
rPAD/2948 PAD:8154 PAD:13862 1.5
rPAD/2949 PAD:8151 PAD:8154 0.0751765
rPAD/2950 PAD:8151 PAD:13859 1.5
rPAD/2951 PAD:8149 PAD:13853 0.0751765
rPAD/2952 PAD:8149 PAD:13859 0.0375882
rPAD/2953 PAD:8149 PAD:13857 1.5
rPAD/2954 PAD:8148 PAD:8151 0.0375882
rPAD/2955 PAD:8148 PAD:8149 1.5
rPAD/2956 PAD:8145 PAD:8148 0.0751765
rPAD/2957 PAD:8145 PAD:13853 1.5
rPAD/2958 PAD:8142 PAD:8145 0.0375882
rPAD/2959 PAD:8142 PAD:13850 1.5
rPAD/2960 PAD:8140 PAD:13850 0.0751765
rPAD/2961 PAD:8140 PAD:13848 1.5
rPAD/2962 PAD:8139 PAD:8142 0.0751765
rPAD/2963 PAD:8139 PAD:8140 1.5
rPAD/2964 PAD:8137 PAD:8140 0.0375882
rPAD/2965 PAD:8137 PAD:13845 1.5
rPAD/2966 PAD:8136 PAD:8139 0.0375882
rPAD/2967 PAD:8136 PAD:8137 1.5
rPAD/2968 PAD:8134 PAD:8137 0.0751765
rPAD/2969 PAD:8134 PAD:13842 1.5
rPAD/2970 PAD:8133 PAD:8136 0.0751765
rPAD/2971 PAD:8133 PAD:8134 1.5
rPAD/2972 PAD:8131 PAD:8134 0.0375882
rPAD/2973 PAD:8131 PAD:13839 1.5
rPAD/2974 PAD:8130 PAD:8133 0.0375882
rPAD/2975 PAD:8130 PAD:8131 1.5
rPAD/2976 PAD:8128 PAD:8131 0.0751765
rPAD/2977 PAD:8128 PAD:13836 1.5
rPAD/2978 PAD:8127 PAD:8130 0.0751765
rPAD/2979 PAD:8127 PAD:8128 1.5
rPAD/2980 PAD:8125 PAD:13829 0.0751765
rPAD/2981 PAD:8125 PAD:8128 0.0375882
rPAD/2982 PAD:8125 PAD:13833 1.5
rPAD/2983 PAD:8124 PAD:8127 0.0375882
rPAD/2984 PAD:8124 PAD:8125 1.5
rPAD/2985 PAD:8121 PAD:8124 0.0751765
rPAD/2986 PAD:8121 PAD:13829 1.5
rPAD/2987 PAD:8119 PAD:13829 0.0375882
rPAD/2988 PAD:8119 PAD:13827 1.5
rPAD/2989 PAD:8118 PAD:8121 0.0375882
rPAD/2990 PAD:8118 PAD:8119 1.5
rPAD/2991 PAD:8116 PAD:8119 0.0751765
rPAD/2992 PAD:8116 PAD:13824 1.5
rPAD/2993 PAD:8115 PAD:8118 0.0751765
rPAD/2994 PAD:8115 PAD:8116 1.5
rPAD/2995 PAD:8113 PAD:13817 0.0751765
rPAD/2996 PAD:8113 PAD:8116 0.0375882
rPAD/2997 PAD:8113 PAD:13821 1.5
rPAD/2998 PAD:8112 PAD:8115 0.0375882
rPAD/2999 PAD:8112 PAD:8113 1.5
rPAD/3000 PAD:8109 PAD:8112 0.0751765
rPAD/3001 PAD:8109 PAD:13817 1.5
rPAD/3002 PAD:8106 PAD:8109 0.0375882
rPAD/3003 PAD:8106 PAD:13814 1.5
rPAD/3004 PAD:8103 PAD:8106 0.0751765
rPAD/3005 PAD:8103 PAD:13811 1.5
rPAD/3006 PAD:8100 PAD:8103 0.0375882
rPAD/3007 PAD:8100 PAD:13808 1.5
rPAD/3008 PAD:8097 PAD:8100 0.0751765
rPAD/3009 PAD:8097 PAD:13805 1.5
rPAD/3010 PAD:8095 PAD:13805 0.0375882
rPAD/3011 PAD:8095 PAD:13803 1.5
rPAD/3012 PAD:8094 PAD:8097 0.0375882
rPAD/3013 PAD:8094 PAD:8095 1.5
rPAD/3014 PAD:8092 PAD:13796 0.0375882
rPAD/3015 PAD:8092 PAD:8095 0.0751765
rPAD/3016 PAD:8092 PAD:13800 1.5
rPAD/3017 PAD:8091 PAD:8094 0.0751765
rPAD/3018 PAD:8091 PAD:8092 1.5
rPAD/3019 PAD:8088 PAD:8091 0.0375882
rPAD/3020 PAD:8088 PAD:13796 1.5
rPAD/3021 PAD:8086 PAD:13796 0.0751765
rPAD/3022 PAD:8086 PAD:13794 1.5
rPAD/3023 PAD:8085 PAD:8088 0.0751765
rPAD/3024 PAD:8085 PAD:8086 1.5
rPAD/3025 PAD:8083 PAD:8086 0.0375882
rPAD/3026 PAD:8083 PAD:13791 1.5
rPAD/3027 PAD:8082 PAD:8085 0.0375882
rPAD/3028 PAD:8082 PAD:8083 1.5
rPAD/3029 PAD:8080 PAD:8083 0.0751765
rPAD/3030 PAD:8080 PAD:13788 1.5
rPAD/3031 PAD:8079 PAD:8082 0.0751765
rPAD/3032 PAD:8079 PAD:8080 1.5
rPAD/3033 PAD:8077 PAD:8080 0.0375882
rPAD/3034 PAD:8077 PAD:13785 1.5
rPAD/3035 PAD:8076 PAD:8079 0.0375882
rPAD/3036 PAD:8076 PAD:8077 1.5
rPAD/3037 PAD:8074 PAD:8077 0.0751765
rPAD/3038 PAD:8074 PAD:13782 1.5
rPAD/3039 PAD:8073 PAD:8076 0.0751765
rPAD/3040 PAD:8073 PAD:8074 1.5
rPAD/3041 PAD:8071 PAD:13775 0.0751765
rPAD/3042 PAD:8071 PAD:8074 0.0375882
rPAD/3043 PAD:8071 PAD:13779 1.5
rPAD/3044 PAD:8070 PAD:8073 0.0375882
rPAD/3045 PAD:8070 PAD:8071 1.5
rPAD/3046 PAD:8067 PAD:8070 0.0751765
rPAD/3047 PAD:8067 PAD:13775 1.5
rPAD/3048 PAD:8065 PAD:13775 0.0375882
rPAD/3049 PAD:8065 PAD:13773 1.5
rPAD/3050 PAD:8064 PAD:8067 0.0375882
rPAD/3051 PAD:8064 PAD:8065 1.5
rPAD/3052 PAD:8062 PAD:8065 0.0751765
rPAD/3053 PAD:8062 PAD:13770 1.5
rPAD/3054 PAD:8061 PAD:8064 0.0751765
rPAD/3055 PAD:8061 PAD:8062 1.5
rPAD/3056 PAD:8059 PAD:8062 0.0375882
rPAD/3057 PAD:8059 PAD:13767 1.5
rPAD/3058 PAD:8058 PAD:8061 0.0375882
rPAD/3059 PAD:8058 PAD:8059 1.5
rPAD/3060 PAD:8056 PAD:8059 0.0751765
rPAD/3061 PAD:8056 PAD:13764 1.5
rPAD/3062 PAD:8055 PAD:8058 0.0751765
rPAD/3063 PAD:8055 PAD:8056 1.5
rPAD/3064 PAD:8053 PAD:8056 0.0375882
rPAD/3065 PAD:8053 PAD:13761 1.5
rPAD/3066 PAD:8052 PAD:8055 0.0375882
rPAD/3067 PAD:8052 PAD:8053 1.5
rPAD/3068 PAD:8050 PAD:8053 0.0751765
rPAD/3069 PAD:8050 PAD:13758 1.5
rPAD/3070 PAD:8049 PAD:8052 0.0751765
rPAD/3071 PAD:8049 PAD:8050 1.5
rPAD/3072 PAD:8047 PAD:8050 0.0375882
rPAD/3073 PAD:8047 PAD:13755 1.5
rPAD/3074 PAD:8046 PAD:8049 0.0375882
rPAD/3075 PAD:8046 PAD:8047 1.5
rPAD/3076 PAD:8044 PAD:14966 0.0283817
rPAD/3077 PAD:8044 PAD:8047 0.0751765
rPAD/3078 PAD:8044 PAD:13752 1.5
rPAD/3079 PAD:8043 PAD:9263 0.0378785
rPAD/3080 PAD:8043 PAD:8046 0.0751765
rPAD/3081 PAD:8043 PAD:8044 1.5
rPAD/3082 PAD:8039 PAD:13579 0.0100588
rPAD/3083 PAD:8039 PAD:13747 1.5
rPAD/3084 PAD:8038 PAD:9418 0.0670908
rPAD/3085 PAD:8038 PAD:8039 1.5
rPAD/3086 PAD:8036 PAD:8039 0.0751765
rPAD/3087 PAD:8036 PAD:13744 1.5
rPAD/3088 PAD:8035 PAD:8038 0.0751765
rPAD/3089 PAD:8035 PAD:8036 1.5
rPAD/3090 PAD:8033 PAD:13737 0.0751765
rPAD/3091 PAD:8033 PAD:8036 0.0375882
rPAD/3092 PAD:8033 PAD:13741 1.5
rPAD/3093 PAD:8032 PAD:8035 0.0375882
rPAD/3094 PAD:8032 PAD:8033 1.5
rPAD/3095 PAD:8029 PAD:8032 0.0751765
rPAD/3096 PAD:8029 PAD:13737 1.5
rPAD/3097 PAD:8027 PAD:13737 0.0375882
rPAD/3098 PAD:8027 PAD:13735 1.5
rPAD/3099 PAD:8026 PAD:8029 0.0375882
rPAD/3100 PAD:8026 PAD:8027 1.5
rPAD/3101 PAD:8024 PAD:8027 0.0751765
rPAD/3102 PAD:8024 PAD:13732 1.5
rPAD/3103 PAD:8023 PAD:8026 0.0751765
rPAD/3104 PAD:8023 PAD:8024 1.5
rPAD/3105 PAD:8021 PAD:8024 0.0375882
rPAD/3106 PAD:8021 PAD:13729 1.5
rPAD/3107 PAD:8020 PAD:8023 0.0375882
rPAD/3108 PAD:8020 PAD:8021 1.5
rPAD/3109 PAD:8018 PAD:8021 0.0751765
rPAD/3110 PAD:8018 PAD:13726 1.5
rPAD/3111 PAD:8017 PAD:8020 0.0751765
rPAD/3112 PAD:8017 PAD:8018 1.5
rPAD/3113 PAD:8015 PAD:8018 0.0375882
rPAD/3114 PAD:8015 PAD:13723 1.5
rPAD/3115 PAD:8014 PAD:8017 0.0375882
rPAD/3116 PAD:8014 PAD:8015 1.5
rPAD/3117 PAD:8012 PAD:8015 0.0751765
rPAD/3118 PAD:8012 PAD:13720 1.5
rPAD/3119 PAD:8011 PAD:8014 0.0751765
rPAD/3120 PAD:8011 PAD:8012 1.5
rPAD/3121 PAD:8009 PAD:8012 0.0375882
rPAD/3122 PAD:8009 PAD:13717 1.5
rPAD/3123 PAD:8008 PAD:8011 0.0375882
rPAD/3124 PAD:8008 PAD:8009 1.5
rPAD/3125 PAD:8006 PAD:8009 0.0751765
rPAD/3126 PAD:8006 PAD:13714 1.5
rPAD/3127 PAD:8005 PAD:8008 0.0751765
rPAD/3128 PAD:8005 PAD:8006 1.5
rPAD/3129 PAD:8003 PAD:8006 0.0375882
rPAD/3130 PAD:8003 PAD:13711 1.5
rPAD/3131 PAD:8002 PAD:8005 0.0375882
rPAD/3132 PAD:8002 PAD:8003 1.5
rPAD/3133 PAD:8000 PAD:8003 0.0751765
rPAD/3134 PAD:8000 PAD:13708 1.5
rPAD/3135 PAD:7999 PAD:8002 0.0751765
rPAD/3136 PAD:7999 PAD:8000 1.5
rPAD/3137 PAD:7997 PAD:13701 0.0751765
rPAD/3138 PAD:7997 PAD:8000 0.0375882
rPAD/3139 PAD:7997 PAD:13705 1.5
rPAD/3140 PAD:7996 PAD:7999 0.0375882
rPAD/3141 PAD:7996 PAD:7997 1.5
rPAD/3142 PAD:7993 PAD:7996 0.0751765
rPAD/3143 PAD:7993 PAD:13701 1.5
rPAD/3144 PAD:7991 PAD:13695 0.0751765
rPAD/3145 PAD:7991 PAD:13701 0.0375882
rPAD/3146 PAD:7991 PAD:13699 1.5
rPAD/3147 PAD:7990 PAD:7993 0.0375882
rPAD/3148 PAD:7990 PAD:7991 1.5
rPAD/3149 PAD:7987 PAD:7990 0.0751765
rPAD/3150 PAD:7987 PAD:13695 1.5
rPAD/3151 PAD:7984 PAD:7987 0.0375882
rPAD/3152 PAD:7984 PAD:13692 1.5
rPAD/3153 PAD:7981 PAD:7984 0.0751765
rPAD/3154 PAD:7981 PAD:13689 1.5
rPAD/3155 PAD:7979 PAD:13683 0.0751765
rPAD/3156 PAD:7979 PAD:13689 0.0375882
rPAD/3157 PAD:7979 PAD:13687 1.5
rPAD/3158 PAD:7978 PAD:7981 0.0375882
rPAD/3159 PAD:7978 PAD:7979 1.5
rPAD/3160 PAD:7975 PAD:7978 0.0751765
rPAD/3161 PAD:7975 PAD:13683 1.5
rPAD/3162 PAD:7972 PAD:7975 0.0375882
rPAD/3163 PAD:7972 PAD:13680 1.5
rPAD/3164 PAD:7970 PAD:13680 0.0751765
rPAD/3165 PAD:7970 PAD:13678 1.5
rPAD/3166 PAD:7969 PAD:7972 0.0751765
rPAD/3167 PAD:7969 PAD:7970 1.5
rPAD/3168 PAD:7967 PAD:7970 0.0375882
rPAD/3169 PAD:7967 PAD:13675 1.5
rPAD/3170 PAD:7966 PAD:7969 0.0375882
rPAD/3171 PAD:7966 PAD:7967 1.5
rPAD/3172 PAD:7964 PAD:7967 0.0751765
rPAD/3173 PAD:7964 PAD:13672 1.5
rPAD/3174 PAD:7963 PAD:7966 0.0751765
rPAD/3175 PAD:7963 PAD:7964 1.5
rPAD/3176 PAD:7961 PAD:7964 0.0375882
rPAD/3177 PAD:7961 PAD:13669 1.5
rPAD/3178 PAD:7960 PAD:7963 0.0375882
rPAD/3179 PAD:7960 PAD:7961 1.5
rPAD/3180 PAD:7958 PAD:7961 0.0751765
rPAD/3181 PAD:7958 PAD:13666 1.5
rPAD/3182 PAD:7957 PAD:7960 0.0751765
rPAD/3183 PAD:7957 PAD:7958 1.5
rPAD/3184 PAD:7955 PAD:13659 0.0751765
rPAD/3185 PAD:7955 PAD:7958 0.0375882
rPAD/3186 PAD:7955 PAD:13663 1.5
rPAD/3187 PAD:7954 PAD:7957 0.0375882
rPAD/3188 PAD:7954 PAD:7955 1.5
rPAD/3189 PAD:7951 PAD:7954 0.0751765
rPAD/3190 PAD:7951 PAD:13659 1.5
rPAD/3191 PAD:7949 PAD:13659 0.0375882
rPAD/3192 PAD:7949 PAD:13657 1.5
rPAD/3193 PAD:7948 PAD:7951 0.0375882
rPAD/3194 PAD:7948 PAD:7949 1.5
rPAD/3195 PAD:7946 PAD:7949 0.0751765
rPAD/3196 PAD:7946 PAD:13654 1.5
rPAD/3197 PAD:7945 PAD:7948 0.0751765
rPAD/3198 PAD:7945 PAD:7946 1.5
rPAD/3199 PAD:7943 PAD:13647 0.0751765
rPAD/3200 PAD:7943 PAD:7946 0.0375882
rPAD/3201 PAD:7943 PAD:13651 1.5
rPAD/3202 PAD:7942 PAD:7945 0.0375882
rPAD/3203 PAD:7942 PAD:7943 1.5
rPAD/3204 PAD:7939 PAD:7942 0.0751765
rPAD/3205 PAD:7939 PAD:13647 1.5
rPAD/3206 PAD:7936 PAD:7939 0.0375882
rPAD/3207 PAD:7936 PAD:13644 1.5
rPAD/3208 PAD:7933 PAD:7936 0.0751765
rPAD/3209 PAD:7933 PAD:13641 1.5
rPAD/3210 PAD:7930 PAD:7933 0.0375882
rPAD/3211 PAD:7930 PAD:13638 1.5
rPAD/3212 PAD:7927 PAD:7930 0.0751765
rPAD/3213 PAD:7927 PAD:13635 1.5
rPAD/3214 PAD:7925 PAD:13635 0.0375882
rPAD/3215 PAD:7925 PAD:13633 1.5
rPAD/3216 PAD:7924 PAD:7927 0.0375882
rPAD/3217 PAD:7924 PAD:7925 1.5
rPAD/3218 PAD:7922 PAD:13626 0.0375882
rPAD/3219 PAD:7922 PAD:7925 0.0751765
rPAD/3220 PAD:7922 PAD:13630 1.5
rPAD/3221 PAD:7921 PAD:7924 0.0751765
rPAD/3222 PAD:7921 PAD:7922 1.5
rPAD/3223 PAD:7918 PAD:7921 0.0375882
rPAD/3224 PAD:7918 PAD:13626 1.5
rPAD/3225 PAD:7916 PAD:13626 0.0751765
rPAD/3226 PAD:7916 PAD:13624 1.5
rPAD/3227 PAD:7915 PAD:7918 0.0751765
rPAD/3228 PAD:7915 PAD:7916 1.5
rPAD/3229 PAD:7913 PAD:7916 0.0375882
rPAD/3230 PAD:7913 PAD:13621 1.5
rPAD/3231 PAD:7912 PAD:7915 0.0375882
rPAD/3232 PAD:7912 PAD:7913 1.5
rPAD/3233 PAD:7910 PAD:7913 0.0751765
rPAD/3234 PAD:7910 PAD:13618 1.5
rPAD/3235 PAD:7909 PAD:7912 0.0751765
rPAD/3236 PAD:7909 PAD:7910 1.5
rPAD/3237 PAD:7907 PAD:7910 0.0375882
rPAD/3238 PAD:7907 PAD:13615 1.5
rPAD/3239 PAD:7906 PAD:7909 0.0375882
rPAD/3240 PAD:7906 PAD:7907 1.5
rPAD/3241 PAD:7904 PAD:7907 0.0751765
rPAD/3242 PAD:7904 PAD:13612 1.5
rPAD/3243 PAD:7903 PAD:7906 0.0751765
rPAD/3244 PAD:7903 PAD:7904 1.5
rPAD/3245 PAD:7901 PAD:13605 0.0751765
rPAD/3246 PAD:7901 PAD:7904 0.0375882
rPAD/3247 PAD:7901 PAD:13609 1.5
rPAD/3248 PAD:7900 PAD:7903 0.0375882
rPAD/3249 PAD:7900 PAD:7901 1.5
rPAD/3250 PAD:7897 PAD:7900 0.0751765
rPAD/3251 PAD:7897 PAD:13605 1.5
rPAD/3252 PAD:7895 PAD:13605 0.0375882
rPAD/3253 PAD:7895 PAD:13603 1.5
rPAD/3254 PAD:7894 PAD:7897 0.0375882
rPAD/3255 PAD:7894 PAD:7895 1.5
rPAD/3256 PAD:7892 PAD:7895 0.0751765
rPAD/3257 PAD:7892 PAD:13600 1.5
rPAD/3258 PAD:7891 PAD:7894 0.0751765
rPAD/3259 PAD:7891 PAD:7892 1.5
rPAD/3260 PAD:7889 PAD:7892 0.0375882
rPAD/3261 PAD:7889 PAD:13597 1.5
rPAD/3262 PAD:7888 PAD:7891 0.0375882
rPAD/3263 PAD:7888 PAD:7889 1.5
rPAD/3264 PAD:7886 PAD:7889 0.0751765
rPAD/3265 PAD:7886 PAD:13594 1.5
rPAD/3266 PAD:7885 PAD:7888 0.0751765
rPAD/3267 PAD:7885 PAD:7886 1.5
rPAD/3268 PAD:7883 PAD:7886 0.0375882
rPAD/3269 PAD:7883 PAD:13591 1.5
rPAD/3270 PAD:7882 PAD:7885 0.0375882
rPAD/3271 PAD:7882 PAD:7883 1.5
rPAD/3272 PAD:7880 PAD:7883 0.0751765
rPAD/3273 PAD:7880 PAD:13588 1.5
rPAD/3274 PAD:7879 PAD:7882 0.0751765
rPAD/3275 PAD:7879 PAD:7880 1.5
rPAD/3276 PAD:7877 PAD:7880 0.0375882
rPAD/3277 PAD:7877 PAD:13585 1.5
rPAD/3278 PAD:7876 PAD:7879 0.0375882
rPAD/3279 PAD:7876 PAD:7877 1.5
rPAD/3280 PAD:7874 PAD:14961 0.0283817
rPAD/3281 PAD:7874 PAD:7877 0.0751765
rPAD/3282 PAD:7874 PAD:13582 1.5
rPAD/3283 PAD:7873 PAD:9256 0.0378785
rPAD/3284 PAD:7873 PAD:7876 0.0751765
rPAD/3285 PAD:7873 PAD:7874 1.5
rPAD/3286 PAD:7869 PAD:13409 0.0100588
rPAD/3287 PAD:7869 PAD:13577 1.5
rPAD/3288 PAD:7868 PAD:9414 0.0670908
rPAD/3289 PAD:7868 PAD:7869 1.5
rPAD/3290 PAD:7866 PAD:7869 0.0751765
rPAD/3291 PAD:7866 PAD:13574 1.5
rPAD/3292 PAD:7865 PAD:7868 0.0751765
rPAD/3293 PAD:7865 PAD:7866 1.5
rPAD/3294 PAD:7863 PAD:13567 0.0751765
rPAD/3295 PAD:7863 PAD:7866 0.0375882
rPAD/3296 PAD:7863 PAD:13571 1.5
rPAD/3297 PAD:7862 PAD:7865 0.0375882
rPAD/3298 PAD:7862 PAD:7863 1.5
rPAD/3299 PAD:7859 PAD:7862 0.0751765
rPAD/3300 PAD:7859 PAD:13567 1.5
rPAD/3301 PAD:7857 PAD:13567 0.0375882
rPAD/3302 PAD:7857 PAD:13565 1.5
rPAD/3303 PAD:7856 PAD:7859 0.0375882
rPAD/3304 PAD:7856 PAD:7857 1.5
rPAD/3305 PAD:7854 PAD:7857 0.0751765
rPAD/3306 PAD:7854 PAD:13562 1.5
rPAD/3307 PAD:7853 PAD:7856 0.0751765
rPAD/3308 PAD:7853 PAD:7854 1.5
rPAD/3309 PAD:7851 PAD:7854 0.0375882
rPAD/3310 PAD:7851 PAD:13559 1.5
rPAD/3311 PAD:7850 PAD:7853 0.0375882
rPAD/3312 PAD:7850 PAD:7851 1.5
rPAD/3313 PAD:7848 PAD:7851 0.0751765
rPAD/3314 PAD:7848 PAD:13556 1.5
rPAD/3315 PAD:7847 PAD:7850 0.0751765
rPAD/3316 PAD:7847 PAD:7848 1.5
rPAD/3317 PAD:7845 PAD:7848 0.0375882
rPAD/3318 PAD:7845 PAD:13553 1.5
rPAD/3319 PAD:7844 PAD:7847 0.0375882
rPAD/3320 PAD:7844 PAD:7845 1.5
rPAD/3321 PAD:7842 PAD:7845 0.0751765
rPAD/3322 PAD:7842 PAD:13550 1.5
rPAD/3323 PAD:7841 PAD:7844 0.0751765
rPAD/3324 PAD:7841 PAD:7842 1.5
rPAD/3325 PAD:7839 PAD:7842 0.0375882
rPAD/3326 PAD:7839 PAD:13547 1.5
rPAD/3327 PAD:7838 PAD:7841 0.0375882
rPAD/3328 PAD:7838 PAD:7839 1.5
rPAD/3329 PAD:7836 PAD:7839 0.0751765
rPAD/3330 PAD:7836 PAD:13544 1.5
rPAD/3331 PAD:7835 PAD:7838 0.0751765
rPAD/3332 PAD:7835 PAD:7836 1.5
rPAD/3333 PAD:7833 PAD:7836 0.0375882
rPAD/3334 PAD:7833 PAD:13541 1.5
rPAD/3335 PAD:7832 PAD:7835 0.0375882
rPAD/3336 PAD:7832 PAD:7833 1.5
rPAD/3337 PAD:7830 PAD:7833 0.0751765
rPAD/3338 PAD:7830 PAD:13538 1.5
rPAD/3339 PAD:7829 PAD:7832 0.0751765
rPAD/3340 PAD:7829 PAD:7830 1.5
rPAD/3341 PAD:7827 PAD:13531 0.0751765
rPAD/3342 PAD:7827 PAD:7830 0.0375882
rPAD/3343 PAD:7827 PAD:13535 1.5
rPAD/3344 PAD:7826 PAD:7829 0.0375882
rPAD/3345 PAD:7826 PAD:7827 1.5
rPAD/3346 PAD:7823 PAD:7826 0.0751765
rPAD/3347 PAD:7823 PAD:13531 1.5
rPAD/3348 PAD:7821 PAD:13525 0.0751765
rPAD/3349 PAD:7821 PAD:13531 0.0375882
rPAD/3350 PAD:7821 PAD:13529 1.5
rPAD/3351 PAD:7820 PAD:7823 0.0375882
rPAD/3352 PAD:7820 PAD:7821 1.5
rPAD/3353 PAD:7817 PAD:7820 0.0751765
rPAD/3354 PAD:7817 PAD:13525 1.5
rPAD/3355 PAD:7814 PAD:7817 0.0375882
rPAD/3356 PAD:7814 PAD:13522 1.5
rPAD/3357 PAD:7811 PAD:7814 0.0751765
rPAD/3358 PAD:7811 PAD:13519 1.5
rPAD/3359 PAD:7809 PAD:13513 0.0751765
rPAD/3360 PAD:7809 PAD:13519 0.0375882
rPAD/3361 PAD:7809 PAD:13517 1.5
rPAD/3362 PAD:7808 PAD:7811 0.0375882
rPAD/3363 PAD:7808 PAD:7809 1.5
rPAD/3364 PAD:7805 PAD:7808 0.0751765
rPAD/3365 PAD:7805 PAD:13513 1.5
rPAD/3366 PAD:7802 PAD:7805 0.0375882
rPAD/3367 PAD:7802 PAD:13510 1.5
rPAD/3368 PAD:7800 PAD:13510 0.0751765
rPAD/3369 PAD:7800 PAD:13508 1.5
rPAD/3370 PAD:7799 PAD:7802 0.0751765
rPAD/3371 PAD:7799 PAD:7800 1.5
rPAD/3372 PAD:7797 PAD:7800 0.0375882
rPAD/3373 PAD:7797 PAD:13505 1.5
rPAD/3374 PAD:7796 PAD:7799 0.0375882
rPAD/3375 PAD:7796 PAD:7797 1.5
rPAD/3376 PAD:7794 PAD:7797 0.0751765
rPAD/3377 PAD:7794 PAD:13502 1.5
rPAD/3378 PAD:7793 PAD:7796 0.0751765
rPAD/3379 PAD:7793 PAD:7794 1.5
rPAD/3380 PAD:7791 PAD:7794 0.0375882
rPAD/3381 PAD:7791 PAD:13499 1.5
rPAD/3382 PAD:7790 PAD:7793 0.0375882
rPAD/3383 PAD:7790 PAD:7791 1.5
rPAD/3384 PAD:7788 PAD:7791 0.0751765
rPAD/3385 PAD:7788 PAD:13496 1.5
rPAD/3386 PAD:7787 PAD:7790 0.0751765
rPAD/3387 PAD:7787 PAD:7788 1.5
rPAD/3388 PAD:7785 PAD:13489 0.0751765
rPAD/3389 PAD:7785 PAD:7788 0.0375882
rPAD/3390 PAD:7785 PAD:13493 1.5
rPAD/3391 PAD:7784 PAD:7787 0.0375882
rPAD/3392 PAD:7784 PAD:7785 1.5
rPAD/3393 PAD:7781 PAD:7784 0.0751765
rPAD/3394 PAD:7781 PAD:13489 1.5
rPAD/3395 PAD:7779 PAD:13489 0.0375882
rPAD/3396 PAD:7779 PAD:13487 1.5
rPAD/3397 PAD:7778 PAD:7781 0.0375882
rPAD/3398 PAD:7778 PAD:7779 1.5
rPAD/3399 PAD:7776 PAD:7779 0.0751765
rPAD/3400 PAD:7776 PAD:13484 1.5
rPAD/3401 PAD:7775 PAD:7778 0.0751765
rPAD/3402 PAD:7775 PAD:7776 1.5
rPAD/3403 PAD:7773 PAD:13477 0.0751765
rPAD/3404 PAD:7773 PAD:7776 0.0375882
rPAD/3405 PAD:7773 PAD:13481 1.5
rPAD/3406 PAD:7772 PAD:7775 0.0375882
rPAD/3407 PAD:7772 PAD:7773 1.5
rPAD/3408 PAD:7769 PAD:7772 0.0751765
rPAD/3409 PAD:7769 PAD:13477 1.5
rPAD/3410 PAD:7766 PAD:7769 0.0375882
rPAD/3411 PAD:7766 PAD:13474 1.5
rPAD/3412 PAD:7763 PAD:7766 0.0751765
rPAD/3413 PAD:7763 PAD:13471 1.5
rPAD/3414 PAD:7760 PAD:7763 0.0375882
rPAD/3415 PAD:7760 PAD:13468 1.5
rPAD/3416 PAD:7757 PAD:7760 0.0751765
rPAD/3417 PAD:7757 PAD:13465 1.5
rPAD/3418 PAD:7755 PAD:13465 0.0375882
rPAD/3419 PAD:7755 PAD:13463 1.5
rPAD/3420 PAD:7754 PAD:7757 0.0375882
rPAD/3421 PAD:7754 PAD:7755 1.5
rPAD/3422 PAD:7752 PAD:13456 0.0375882
rPAD/3423 PAD:7752 PAD:7755 0.0751765
rPAD/3424 PAD:7752 PAD:13460 1.5
rPAD/3425 PAD:7751 PAD:7754 0.0751765
rPAD/3426 PAD:7751 PAD:7752 1.5
rPAD/3427 PAD:7748 PAD:7751 0.0375882
rPAD/3428 PAD:7748 PAD:13456 1.5
rPAD/3429 PAD:7746 PAD:13456 0.0751765
rPAD/3430 PAD:7746 PAD:13454 1.5
rPAD/3431 PAD:7745 PAD:7748 0.0751765
rPAD/3432 PAD:7745 PAD:7746 1.5
rPAD/3433 PAD:7743 PAD:7746 0.0375882
rPAD/3434 PAD:7743 PAD:13451 1.5
rPAD/3435 PAD:7742 PAD:7745 0.0375882
rPAD/3436 PAD:7742 PAD:7743 1.5
rPAD/3437 PAD:7740 PAD:7743 0.0751765
rPAD/3438 PAD:7740 PAD:13448 1.5
rPAD/3439 PAD:7739 PAD:7742 0.0751765
rPAD/3440 PAD:7739 PAD:7740 1.5
rPAD/3441 PAD:7737 PAD:7740 0.0375882
rPAD/3442 PAD:7737 PAD:13445 1.5
rPAD/3443 PAD:7736 PAD:7739 0.0375882
rPAD/3444 PAD:7736 PAD:7737 1.5
rPAD/3445 PAD:7734 PAD:7737 0.0751765
rPAD/3446 PAD:7734 PAD:13442 1.5
rPAD/3447 PAD:7733 PAD:7736 0.0751765
rPAD/3448 PAD:7733 PAD:7734 1.5
rPAD/3449 PAD:7731 PAD:13435 0.0751765
rPAD/3450 PAD:7731 PAD:7734 0.0375882
rPAD/3451 PAD:7731 PAD:13439 1.5
rPAD/3452 PAD:7730 PAD:7733 0.0375882
rPAD/3453 PAD:7730 PAD:7731 1.5
rPAD/3454 PAD:7727 PAD:7730 0.0751765
rPAD/3455 PAD:7727 PAD:13435 1.5
rPAD/3456 PAD:7725 PAD:13435 0.0375882
rPAD/3457 PAD:7725 PAD:13433 1.5
rPAD/3458 PAD:7724 PAD:7727 0.0375882
rPAD/3459 PAD:7724 PAD:7725 1.5
rPAD/3460 PAD:7722 PAD:7725 0.0751765
rPAD/3461 PAD:7722 PAD:13430 1.5
rPAD/3462 PAD:7721 PAD:7724 0.0751765
rPAD/3463 PAD:7721 PAD:7722 1.5
rPAD/3464 PAD:7719 PAD:7722 0.0375882
rPAD/3465 PAD:7719 PAD:13427 1.5
rPAD/3466 PAD:7718 PAD:7721 0.0375882
rPAD/3467 PAD:7718 PAD:7719 1.5
rPAD/3468 PAD:7716 PAD:7719 0.0751765
rPAD/3469 PAD:7716 PAD:13424 1.5
rPAD/3470 PAD:7715 PAD:7718 0.0751765
rPAD/3471 PAD:7715 PAD:7716 1.5
rPAD/3472 PAD:7713 PAD:7716 0.0375882
rPAD/3473 PAD:7713 PAD:13421 1.5
rPAD/3474 PAD:7712 PAD:7715 0.0375882
rPAD/3475 PAD:7712 PAD:7713 1.5
rPAD/3476 PAD:7710 PAD:7713 0.0751765
rPAD/3477 PAD:7710 PAD:13418 1.5
rPAD/3478 PAD:7709 PAD:7712 0.0751765
rPAD/3479 PAD:7709 PAD:7710 1.5
rPAD/3480 PAD:7707 PAD:7710 0.0375882
rPAD/3481 PAD:7707 PAD:13415 1.5
rPAD/3482 PAD:7706 PAD:7709 0.0375882
rPAD/3483 PAD:7706 PAD:7707 1.5
rPAD/3484 PAD:7704 PAD:14955 0.0283817
rPAD/3485 PAD:7704 PAD:7707 0.0751765
rPAD/3486 PAD:7704 PAD:13412 1.5
rPAD/3487 PAD:7703 PAD:9249 0.0378785
rPAD/3488 PAD:7703 PAD:7706 0.0751765
rPAD/3489 PAD:7703 PAD:7704 1.5
rPAD/3490 PAD:7699 PAD:13239 0.0100588
rPAD/3491 PAD:7699 PAD:13407 1.5
rPAD/3492 PAD:7698 PAD:9409 0.0670908
rPAD/3493 PAD:7698 PAD:7699 1.5
rPAD/3494 PAD:7696 PAD:7699 0.0751765
rPAD/3495 PAD:7696 PAD:13404 1.5
rPAD/3496 PAD:7695 PAD:7698 0.0751765
rPAD/3497 PAD:7695 PAD:7696 1.5
rPAD/3498 PAD:7693 PAD:13397 0.0751765
rPAD/3499 PAD:7693 PAD:7696 0.0375882
rPAD/3500 PAD:7693 PAD:13401 1.5
rPAD/3501 PAD:7692 PAD:7695 0.0375882
rPAD/3502 PAD:7692 PAD:7693 1.5
rPAD/3503 PAD:7689 PAD:7692 0.0751765
rPAD/3504 PAD:7689 PAD:13397 1.5
rPAD/3505 PAD:7687 PAD:13397 0.0375882
rPAD/3506 PAD:7687 PAD:13395 1.5
rPAD/3507 PAD:7686 PAD:7689 0.0375882
rPAD/3508 PAD:7686 PAD:7687 1.5
rPAD/3509 PAD:7684 PAD:7687 0.0751765
rPAD/3510 PAD:7684 PAD:13392 1.5
rPAD/3511 PAD:7683 PAD:7686 0.0751765
rPAD/3512 PAD:7683 PAD:7684 1.5
rPAD/3513 PAD:7681 PAD:7684 0.0375882
rPAD/3514 PAD:7681 PAD:13389 1.5
rPAD/3515 PAD:7680 PAD:7683 0.0375882
rPAD/3516 PAD:7680 PAD:7681 1.5
rPAD/3517 PAD:7678 PAD:7681 0.0751765
rPAD/3518 PAD:7678 PAD:13386 1.5
rPAD/3519 PAD:7677 PAD:7680 0.0751765
rPAD/3520 PAD:7677 PAD:7678 1.5
rPAD/3521 PAD:7675 PAD:7678 0.0375882
rPAD/3522 PAD:7675 PAD:13383 1.5
rPAD/3523 PAD:7674 PAD:7677 0.0375882
rPAD/3524 PAD:7674 PAD:7675 1.5
rPAD/3525 PAD:7672 PAD:7675 0.0751765
rPAD/3526 PAD:7672 PAD:13380 1.5
rPAD/3527 PAD:7671 PAD:7674 0.0751765
rPAD/3528 PAD:7671 PAD:7672 1.5
rPAD/3529 PAD:7669 PAD:7672 0.0375882
rPAD/3530 PAD:7669 PAD:13377 1.5
rPAD/3531 PAD:7668 PAD:7671 0.0375882
rPAD/3532 PAD:7668 PAD:7669 1.5
rPAD/3533 PAD:7666 PAD:7669 0.0751765
rPAD/3534 PAD:7666 PAD:13374 1.5
rPAD/3535 PAD:7665 PAD:7668 0.0751765
rPAD/3536 PAD:7665 PAD:7666 1.5
rPAD/3537 PAD:7663 PAD:7666 0.0375882
rPAD/3538 PAD:7663 PAD:13371 1.5
rPAD/3539 PAD:7662 PAD:7665 0.0375882
rPAD/3540 PAD:7662 PAD:7663 1.5
rPAD/3541 PAD:7660 PAD:7663 0.0751765
rPAD/3542 PAD:7660 PAD:13368 1.5
rPAD/3543 PAD:7659 PAD:7662 0.0751765
rPAD/3544 PAD:7659 PAD:7660 1.5
rPAD/3545 PAD:7657 PAD:13361 0.0751765
rPAD/3546 PAD:7657 PAD:7660 0.0375882
rPAD/3547 PAD:7657 PAD:13365 1.5
rPAD/3548 PAD:7656 PAD:7659 0.0375882
rPAD/3549 PAD:7656 PAD:7657 1.5
rPAD/3550 PAD:7653 PAD:7656 0.0751765
rPAD/3551 PAD:7653 PAD:13361 1.5
rPAD/3552 PAD:7651 PAD:13355 0.0751765
rPAD/3553 PAD:7651 PAD:13361 0.0375882
rPAD/3554 PAD:7651 PAD:13359 1.5
rPAD/3555 PAD:7650 PAD:7653 0.0375882
rPAD/3556 PAD:7650 PAD:7651 1.5
rPAD/3557 PAD:7647 PAD:7650 0.0751765
rPAD/3558 PAD:7647 PAD:13355 1.5
rPAD/3559 PAD:7644 PAD:7647 0.0375882
rPAD/3560 PAD:7644 PAD:13352 1.5
rPAD/3561 PAD:7641 PAD:7644 0.0751765
rPAD/3562 PAD:7641 PAD:13349 1.5
rPAD/3563 PAD:7639 PAD:13343 0.0751765
rPAD/3564 PAD:7639 PAD:13349 0.0375882
rPAD/3565 PAD:7639 PAD:13347 1.5
rPAD/3566 PAD:7638 PAD:7641 0.0375882
rPAD/3567 PAD:7638 PAD:7639 1.5
rPAD/3568 PAD:7635 PAD:7638 0.0751765
rPAD/3569 PAD:7635 PAD:13343 1.5
rPAD/3570 PAD:7632 PAD:7635 0.0375882
rPAD/3571 PAD:7632 PAD:13340 1.5
rPAD/3572 PAD:7630 PAD:13340 0.0751765
rPAD/3573 PAD:7630 PAD:13338 1.5
rPAD/3574 PAD:7629 PAD:7632 0.0751765
rPAD/3575 PAD:7629 PAD:7630 1.5
rPAD/3576 PAD:7627 PAD:7630 0.0375882
rPAD/3577 PAD:7627 PAD:13335 1.5
rPAD/3578 PAD:7626 PAD:7629 0.0375882
rPAD/3579 PAD:7626 PAD:7627 1.5
rPAD/3580 PAD:7624 PAD:7627 0.0751765
rPAD/3581 PAD:7624 PAD:13332 1.5
rPAD/3582 PAD:7623 PAD:7626 0.0751765
rPAD/3583 PAD:7623 PAD:7624 1.5
rPAD/3584 PAD:7621 PAD:7624 0.0375882
rPAD/3585 PAD:7621 PAD:13329 1.5
rPAD/3586 PAD:7620 PAD:7623 0.0375882
rPAD/3587 PAD:7620 PAD:7621 1.5
rPAD/3588 PAD:7618 PAD:7621 0.0751765
rPAD/3589 PAD:7618 PAD:13326 1.5
rPAD/3590 PAD:7617 PAD:7620 0.0751765
rPAD/3591 PAD:7617 PAD:7618 1.5
rPAD/3592 PAD:7615 PAD:13319 0.0751765
rPAD/3593 PAD:7615 PAD:7618 0.0375882
rPAD/3594 PAD:7615 PAD:13323 1.5
rPAD/3595 PAD:7614 PAD:7617 0.0375882
rPAD/3596 PAD:7614 PAD:7615 1.5
rPAD/3597 PAD:7611 PAD:7614 0.0751765
rPAD/3598 PAD:7611 PAD:13319 1.5
rPAD/3599 PAD:7609 PAD:13319 0.0375882
rPAD/3600 PAD:7609 PAD:13317 1.5
rPAD/3601 PAD:7608 PAD:7611 0.0375882
rPAD/3602 PAD:7608 PAD:7609 1.5
rPAD/3603 PAD:7606 PAD:7609 0.0751765
rPAD/3604 PAD:7606 PAD:13314 1.5
rPAD/3605 PAD:7605 PAD:7608 0.0751765
rPAD/3606 PAD:7605 PAD:7606 1.5
rPAD/3607 PAD:7603 PAD:13307 0.0751765
rPAD/3608 PAD:7603 PAD:7606 0.0375882
rPAD/3609 PAD:7603 PAD:13311 1.5
rPAD/3610 PAD:7602 PAD:7605 0.0375882
rPAD/3611 PAD:7602 PAD:7603 1.5
rPAD/3612 PAD:7599 PAD:7602 0.0751765
rPAD/3613 PAD:7599 PAD:13307 1.5
rPAD/3614 PAD:7596 PAD:7599 0.0375882
rPAD/3615 PAD:7596 PAD:13304 1.5
rPAD/3616 PAD:7593 PAD:7596 0.0751765
rPAD/3617 PAD:7593 PAD:13301 1.5
rPAD/3618 PAD:7590 PAD:7593 0.0375882
rPAD/3619 PAD:7590 PAD:13298 1.5
rPAD/3620 PAD:7587 PAD:7590 0.0751765
rPAD/3621 PAD:7587 PAD:13295 1.5
rPAD/3622 PAD:7585 PAD:13295 0.0375882
rPAD/3623 PAD:7585 PAD:13293 1.5
rPAD/3624 PAD:7584 PAD:7587 0.0375882
rPAD/3625 PAD:7584 PAD:7585 1.5
rPAD/3626 PAD:7582 PAD:13286 0.0375882
rPAD/3627 PAD:7582 PAD:7585 0.0751765
rPAD/3628 PAD:7582 PAD:13290 1.5
rPAD/3629 PAD:7581 PAD:7584 0.0751765
rPAD/3630 PAD:7581 PAD:7582 1.5
rPAD/3631 PAD:7578 PAD:7581 0.0375882
rPAD/3632 PAD:7578 PAD:13286 1.5
rPAD/3633 PAD:7576 PAD:13286 0.0751765
rPAD/3634 PAD:7576 PAD:13284 1.5
rPAD/3635 PAD:7575 PAD:7578 0.0751765
rPAD/3636 PAD:7575 PAD:7576 1.5
rPAD/3637 PAD:7573 PAD:7576 0.0375882
rPAD/3638 PAD:7573 PAD:13281 1.5
rPAD/3639 PAD:7572 PAD:7575 0.0375882
rPAD/3640 PAD:7572 PAD:7573 1.5
rPAD/3641 PAD:7570 PAD:7573 0.0751765
rPAD/3642 PAD:7570 PAD:13278 1.5
rPAD/3643 PAD:7569 PAD:7572 0.0751765
rPAD/3644 PAD:7569 PAD:7570 1.5
rPAD/3645 PAD:7567 PAD:7570 0.0375882
rPAD/3646 PAD:7567 PAD:13275 1.5
rPAD/3647 PAD:7566 PAD:7569 0.0375882
rPAD/3648 PAD:7566 PAD:7567 1.5
rPAD/3649 PAD:7564 PAD:7567 0.0751765
rPAD/3650 PAD:7564 PAD:13272 1.5
rPAD/3651 PAD:7563 PAD:7566 0.0751765
rPAD/3652 PAD:7563 PAD:7564 1.5
rPAD/3653 PAD:7561 PAD:13265 0.0751765
rPAD/3654 PAD:7561 PAD:7564 0.0375882
rPAD/3655 PAD:7561 PAD:13269 1.5
rPAD/3656 PAD:7560 PAD:7563 0.0375882
rPAD/3657 PAD:7560 PAD:7561 1.5
rPAD/3658 PAD:7557 PAD:7560 0.0751765
rPAD/3659 PAD:7557 PAD:13265 1.5
rPAD/3660 PAD:7555 PAD:13265 0.0375882
rPAD/3661 PAD:7555 PAD:13263 1.5
rPAD/3662 PAD:7554 PAD:7557 0.0375882
rPAD/3663 PAD:7554 PAD:7555 1.5
rPAD/3664 PAD:7552 PAD:7555 0.0751765
rPAD/3665 PAD:7552 PAD:13260 1.5
rPAD/3666 PAD:7551 PAD:7554 0.0751765
rPAD/3667 PAD:7551 PAD:7552 1.5
rPAD/3668 PAD:7549 PAD:7552 0.0375882
rPAD/3669 PAD:7549 PAD:13257 1.5
rPAD/3670 PAD:7548 PAD:7551 0.0375882
rPAD/3671 PAD:7548 PAD:7549 1.5
rPAD/3672 PAD:7546 PAD:7549 0.0751765
rPAD/3673 PAD:7546 PAD:13254 1.5
rPAD/3674 PAD:7545 PAD:7548 0.0751765
rPAD/3675 PAD:7545 PAD:7546 1.5
rPAD/3676 PAD:7543 PAD:7546 0.0375882
rPAD/3677 PAD:7543 PAD:13251 1.5
rPAD/3678 PAD:7542 PAD:7545 0.0375882
rPAD/3679 PAD:7542 PAD:7543 1.5
rPAD/3680 PAD:7540 PAD:7543 0.0751765
rPAD/3681 PAD:7540 PAD:13248 1.5
rPAD/3682 PAD:7539 PAD:7542 0.0751765
rPAD/3683 PAD:7539 PAD:7540 1.5
rPAD/3684 PAD:7537 PAD:7540 0.0375882
rPAD/3685 PAD:7537 PAD:13245 1.5
rPAD/3686 PAD:7536 PAD:7539 0.0375882
rPAD/3687 PAD:7536 PAD:7537 1.5
rPAD/3688 PAD:7534 PAD:14949 0.0283817
rPAD/3689 PAD:7534 PAD:7537 0.0751765
rPAD/3690 PAD:7534 PAD:13242 1.5
rPAD/3691 PAD:7533 PAD:9242 0.0378785
rPAD/3692 PAD:7533 PAD:7536 0.0751765
rPAD/3693 PAD:7533 PAD:7534 1.5
rPAD/3694 PAD:7529 PAD:13069 0.0100588
rPAD/3695 PAD:7529 PAD:13237 1.5
rPAD/3696 PAD:7528 PAD:9405 0.0670908
rPAD/3697 PAD:7528 PAD:7529 1.5
rPAD/3698 PAD:7526 PAD:7529 0.0751765
rPAD/3699 PAD:7526 PAD:13234 1.5
rPAD/3700 PAD:7525 PAD:7528 0.0751765
rPAD/3701 PAD:7525 PAD:7526 1.5
rPAD/3702 PAD:7523 PAD:13227 0.0751765
rPAD/3703 PAD:7523 PAD:7526 0.0375882
rPAD/3704 PAD:7523 PAD:13231 1.5
rPAD/3705 PAD:7522 PAD:7525 0.0375882
rPAD/3706 PAD:7522 PAD:7523 1.5
rPAD/3707 PAD:7519 PAD:7522 0.0751765
rPAD/3708 PAD:7519 PAD:13227 1.5
rPAD/3709 PAD:7517 PAD:13227 0.0375882
rPAD/3710 PAD:7517 PAD:13225 1.5
rPAD/3711 PAD:7516 PAD:7519 0.0375882
rPAD/3712 PAD:7516 PAD:7517 1.5
rPAD/3713 PAD:7514 PAD:7517 0.0751765
rPAD/3714 PAD:7514 PAD:13222 1.5
rPAD/3715 PAD:7513 PAD:7516 0.0751765
rPAD/3716 PAD:7513 PAD:7514 1.5
rPAD/3717 PAD:7511 PAD:7514 0.0375882
rPAD/3718 PAD:7511 PAD:13219 1.5
rPAD/3719 PAD:7510 PAD:7513 0.0375882
rPAD/3720 PAD:7510 PAD:7511 1.5
rPAD/3721 PAD:7508 PAD:7511 0.0751765
rPAD/3722 PAD:7508 PAD:13216 1.5
rPAD/3723 PAD:7507 PAD:7510 0.0751765
rPAD/3724 PAD:7507 PAD:7508 1.5
rPAD/3725 PAD:7505 PAD:7508 0.0375882
rPAD/3726 PAD:7505 PAD:13213 1.5
rPAD/3727 PAD:7504 PAD:7507 0.0375882
rPAD/3728 PAD:7504 PAD:7505 1.5
rPAD/3729 PAD:7502 PAD:7505 0.0751765
rPAD/3730 PAD:7502 PAD:13210 1.5
rPAD/3731 PAD:7501 PAD:7504 0.0751765
rPAD/3732 PAD:7501 PAD:7502 1.5
rPAD/3733 PAD:7499 PAD:7502 0.0375882
rPAD/3734 PAD:7499 PAD:13207 1.5
rPAD/3735 PAD:7498 PAD:7501 0.0375882
rPAD/3736 PAD:7498 PAD:7499 1.5
rPAD/3737 PAD:7496 PAD:7499 0.0751765
rPAD/3738 PAD:7496 PAD:13204 1.5
rPAD/3739 PAD:7495 PAD:7498 0.0751765
rPAD/3740 PAD:7495 PAD:7496 1.5
rPAD/3741 PAD:7493 PAD:7496 0.0375882
rPAD/3742 PAD:7493 PAD:13201 1.5
rPAD/3743 PAD:7492 PAD:7495 0.0375882
rPAD/3744 PAD:7492 PAD:7493 1.5
rPAD/3745 PAD:7490 PAD:7493 0.0751765
rPAD/3746 PAD:7490 PAD:13198 1.5
rPAD/3747 PAD:7489 PAD:7492 0.0751765
rPAD/3748 PAD:7489 PAD:7490 1.5
rPAD/3749 PAD:7487 PAD:13191 0.0751765
rPAD/3750 PAD:7487 PAD:7490 0.0375882
rPAD/3751 PAD:7487 PAD:13195 1.5
rPAD/3752 PAD:7486 PAD:7489 0.0375882
rPAD/3753 PAD:7486 PAD:7487 1.5
rPAD/3754 PAD:7483 PAD:7486 0.0751765
rPAD/3755 PAD:7483 PAD:13191 1.5
rPAD/3756 PAD:7481 PAD:13185 0.0751765
rPAD/3757 PAD:7481 PAD:13191 0.0375882
rPAD/3758 PAD:7481 PAD:13189 1.5
rPAD/3759 PAD:7480 PAD:7483 0.0375882
rPAD/3760 PAD:7480 PAD:7481 1.5
rPAD/3761 PAD:7477 PAD:7480 0.0751765
rPAD/3762 PAD:7477 PAD:13185 1.5
rPAD/3763 PAD:7474 PAD:7477 0.0375882
rPAD/3764 PAD:7474 PAD:13182 1.5
rPAD/3765 PAD:7471 PAD:7474 0.0751765
rPAD/3766 PAD:7471 PAD:13179 1.5
rPAD/3767 PAD:7469 PAD:13173 0.0751765
rPAD/3768 PAD:7469 PAD:13179 0.0375882
rPAD/3769 PAD:7469 PAD:13177 1.5
rPAD/3770 PAD:7468 PAD:7471 0.0375882
rPAD/3771 PAD:7468 PAD:7469 1.5
rPAD/3772 PAD:7465 PAD:7468 0.0751765
rPAD/3773 PAD:7465 PAD:13173 1.5
rPAD/3774 PAD:7462 PAD:7465 0.0375882
rPAD/3775 PAD:7462 PAD:13170 1.5
rPAD/3776 PAD:7460 PAD:13170 0.0751765
rPAD/3777 PAD:7460 PAD:13168 1.5
rPAD/3778 PAD:7459 PAD:7462 0.0751765
rPAD/3779 PAD:7459 PAD:7460 1.5
rPAD/3780 PAD:7457 PAD:7460 0.0375882
rPAD/3781 PAD:7457 PAD:13165 1.5
rPAD/3782 PAD:7456 PAD:7459 0.0375882
rPAD/3783 PAD:7456 PAD:7457 1.5
rPAD/3784 PAD:7454 PAD:7457 0.0751765
rPAD/3785 PAD:7454 PAD:13162 1.5
rPAD/3786 PAD:7453 PAD:7456 0.0751765
rPAD/3787 PAD:7453 PAD:7454 1.5
rPAD/3788 PAD:7451 PAD:7454 0.0375882
rPAD/3789 PAD:7451 PAD:13159 1.5
rPAD/3790 PAD:7450 PAD:7453 0.0375882
rPAD/3791 PAD:7450 PAD:7451 1.5
rPAD/3792 PAD:7448 PAD:7451 0.0751765
rPAD/3793 PAD:7448 PAD:13156 1.5
rPAD/3794 PAD:7447 PAD:7450 0.0751765
rPAD/3795 PAD:7447 PAD:7448 1.5
rPAD/3796 PAD:7445 PAD:13149 0.0751765
rPAD/3797 PAD:7445 PAD:7448 0.0375882
rPAD/3798 PAD:7445 PAD:13153 1.5
rPAD/3799 PAD:7444 PAD:7447 0.0375882
rPAD/3800 PAD:7444 PAD:7445 1.5
rPAD/3801 PAD:7441 PAD:7444 0.0751765
rPAD/3802 PAD:7441 PAD:13149 1.5
rPAD/3803 PAD:7439 PAD:13149 0.0375882
rPAD/3804 PAD:7439 PAD:13147 1.5
rPAD/3805 PAD:7438 PAD:7441 0.0375882
rPAD/3806 PAD:7438 PAD:7439 1.5
rPAD/3807 PAD:7436 PAD:7439 0.0751765
rPAD/3808 PAD:7436 PAD:13144 1.5
rPAD/3809 PAD:7435 PAD:7438 0.0751765
rPAD/3810 PAD:7435 PAD:7436 1.5
rPAD/3811 PAD:7433 PAD:13137 0.0751765
rPAD/3812 PAD:7433 PAD:7436 0.0375882
rPAD/3813 PAD:7433 PAD:13141 1.5
rPAD/3814 PAD:7432 PAD:7435 0.0375882
rPAD/3815 PAD:7432 PAD:7433 1.5
rPAD/3816 PAD:7429 PAD:7432 0.0751765
rPAD/3817 PAD:7429 PAD:13137 1.5
rPAD/3818 PAD:7426 PAD:7429 0.0375882
rPAD/3819 PAD:7426 PAD:13134 1.5
rPAD/3820 PAD:7423 PAD:7426 0.0751765
rPAD/3821 PAD:7423 PAD:13131 1.5
rPAD/3822 PAD:7420 PAD:7423 0.0375882
rPAD/3823 PAD:7420 PAD:13128 1.5
rPAD/3824 PAD:7417 PAD:7420 0.0751765
rPAD/3825 PAD:7417 PAD:13125 1.5
rPAD/3826 PAD:7415 PAD:13125 0.0375882
rPAD/3827 PAD:7415 PAD:13123 1.5
rPAD/3828 PAD:7414 PAD:7417 0.0375882
rPAD/3829 PAD:7414 PAD:7415 1.5
rPAD/3830 PAD:7412 PAD:13116 0.0375882
rPAD/3831 PAD:7412 PAD:7415 0.0751765
rPAD/3832 PAD:7412 PAD:13120 1.5
rPAD/3833 PAD:7411 PAD:7414 0.0751765
rPAD/3834 PAD:7411 PAD:7412 1.5
rPAD/3835 PAD:7408 PAD:7411 0.0375882
rPAD/3836 PAD:7408 PAD:13116 1.5
rPAD/3837 PAD:7406 PAD:13116 0.0751765
rPAD/3838 PAD:7406 PAD:13114 1.5
rPAD/3839 PAD:7405 PAD:7408 0.0751765
rPAD/3840 PAD:7405 PAD:7406 1.5
rPAD/3841 PAD:7403 PAD:7406 0.0375882
rPAD/3842 PAD:7403 PAD:13111 1.5
rPAD/3843 PAD:7402 PAD:7405 0.0375882
rPAD/3844 PAD:7402 PAD:7403 1.5
rPAD/3845 PAD:7400 PAD:7403 0.0751765
rPAD/3846 PAD:7400 PAD:13108 1.5
rPAD/3847 PAD:7399 PAD:7402 0.0751765
rPAD/3848 PAD:7399 PAD:7400 1.5
rPAD/3849 PAD:7397 PAD:7400 0.0375882
rPAD/3850 PAD:7397 PAD:13105 1.5
rPAD/3851 PAD:7396 PAD:7399 0.0375882
rPAD/3852 PAD:7396 PAD:7397 1.5
rPAD/3853 PAD:7394 PAD:7397 0.0751765
rPAD/3854 PAD:7394 PAD:13102 1.5
rPAD/3855 PAD:7393 PAD:7396 0.0751765
rPAD/3856 PAD:7393 PAD:7394 1.5
rPAD/3857 PAD:7391 PAD:13095 0.0751765
rPAD/3858 PAD:7391 PAD:7394 0.0375882
rPAD/3859 PAD:7391 PAD:13099 1.5
rPAD/3860 PAD:7390 PAD:7393 0.0375882
rPAD/3861 PAD:7390 PAD:7391 1.5
rPAD/3862 PAD:7387 PAD:7390 0.0751765
rPAD/3863 PAD:7387 PAD:13095 1.5
rPAD/3864 PAD:7385 PAD:13095 0.0375882
rPAD/3865 PAD:7385 PAD:13093 1.5
rPAD/3866 PAD:7384 PAD:7387 0.0375882
rPAD/3867 PAD:7384 PAD:7385 1.5
rPAD/3868 PAD:7382 PAD:7385 0.0751765
rPAD/3869 PAD:7382 PAD:13090 1.5
rPAD/3870 PAD:7381 PAD:7384 0.0751765
rPAD/3871 PAD:7381 PAD:7382 1.5
rPAD/3872 PAD:7379 PAD:7382 0.0375882
rPAD/3873 PAD:7379 PAD:13087 1.5
rPAD/3874 PAD:7378 PAD:7381 0.0375882
rPAD/3875 PAD:7378 PAD:7379 1.5
rPAD/3876 PAD:7376 PAD:7379 0.0751765
rPAD/3877 PAD:7376 PAD:13084 1.5
rPAD/3878 PAD:7375 PAD:7378 0.0751765
rPAD/3879 PAD:7375 PAD:7376 1.5
rPAD/3880 PAD:7373 PAD:7376 0.0375882
rPAD/3881 PAD:7373 PAD:13081 1.5
rPAD/3882 PAD:7372 PAD:7375 0.0375882
rPAD/3883 PAD:7372 PAD:7373 1.5
rPAD/3884 PAD:7370 PAD:7373 0.0751765
rPAD/3885 PAD:7370 PAD:13078 1.5
rPAD/3886 PAD:7369 PAD:7372 0.0751765
rPAD/3887 PAD:7369 PAD:7370 1.5
rPAD/3888 PAD:7367 PAD:7370 0.0375882
rPAD/3889 PAD:7367 PAD:13075 1.5
rPAD/3890 PAD:7366 PAD:7369 0.0375882
rPAD/3891 PAD:7366 PAD:7367 1.5
rPAD/3892 PAD:7364 PAD:14945 0.0283817
rPAD/3893 PAD:7364 PAD:7367 0.0751765
rPAD/3894 PAD:7364 PAD:13072 1.5
rPAD/3895 PAD:7363 PAD:9238 0.0378785
rPAD/3896 PAD:7363 PAD:7366 0.0751765
rPAD/3897 PAD:7363 PAD:7364 1.5
rPAD/3898 PAD:7359 PAD:12899 0.0100588
rPAD/3899 PAD:7359 PAD:13067 1.5
rPAD/3900 PAD:7358 PAD:9401 0.0670908
rPAD/3901 PAD:7358 PAD:7359 1.5
rPAD/3902 PAD:7356 PAD:7359 0.0751765
rPAD/3903 PAD:7356 PAD:13064 1.5
rPAD/3904 PAD:7355 PAD:7358 0.0751765
rPAD/3905 PAD:7355 PAD:7356 1.5
rPAD/3906 PAD:7353 PAD:13057 0.0751765
rPAD/3907 PAD:7353 PAD:7356 0.0375882
rPAD/3908 PAD:7353 PAD:13061 1.5
rPAD/3909 PAD:7352 PAD:7355 0.0375882
rPAD/3910 PAD:7352 PAD:7353 1.5
rPAD/3911 PAD:7349 PAD:7352 0.0751765
rPAD/3912 PAD:7349 PAD:13057 1.5
rPAD/3913 PAD:7347 PAD:13057 0.0375882
rPAD/3914 PAD:7347 PAD:13055 1.5
rPAD/3915 PAD:7346 PAD:7349 0.0375882
rPAD/3916 PAD:7346 PAD:7347 1.5
rPAD/3917 PAD:7344 PAD:7347 0.0751765
rPAD/3918 PAD:7344 PAD:13052 1.5
rPAD/3919 PAD:7343 PAD:7346 0.0751765
rPAD/3920 PAD:7343 PAD:7344 1.5
rPAD/3921 PAD:7341 PAD:7344 0.0375882
rPAD/3922 PAD:7341 PAD:13049 1.5
rPAD/3923 PAD:7340 PAD:7343 0.0375882
rPAD/3924 PAD:7340 PAD:7341 1.5
rPAD/3925 PAD:7338 PAD:7341 0.0751765
rPAD/3926 PAD:7338 PAD:13046 1.5
rPAD/3927 PAD:7337 PAD:7340 0.0751765
rPAD/3928 PAD:7337 PAD:7338 1.5
rPAD/3929 PAD:7335 PAD:7338 0.0375882
rPAD/3930 PAD:7335 PAD:13043 1.5
rPAD/3931 PAD:7334 PAD:7337 0.0375882
rPAD/3932 PAD:7334 PAD:7335 1.5
rPAD/3933 PAD:7332 PAD:7335 0.0751765
rPAD/3934 PAD:7332 PAD:13040 1.5
rPAD/3935 PAD:7331 PAD:7334 0.0751765
rPAD/3936 PAD:7331 PAD:7332 1.5
rPAD/3937 PAD:7329 PAD:7332 0.0375882
rPAD/3938 PAD:7329 PAD:13037 1.5
rPAD/3939 PAD:7328 PAD:7331 0.0375882
rPAD/3940 PAD:7328 PAD:7329 1.5
rPAD/3941 PAD:7326 PAD:7329 0.0751765
rPAD/3942 PAD:7326 PAD:13034 1.5
rPAD/3943 PAD:7325 PAD:7328 0.0751765
rPAD/3944 PAD:7325 PAD:7326 1.5
rPAD/3945 PAD:7323 PAD:7326 0.0375882
rPAD/3946 PAD:7323 PAD:13031 1.5
rPAD/3947 PAD:7322 PAD:7325 0.0375882
rPAD/3948 PAD:7322 PAD:7323 1.5
rPAD/3949 PAD:7320 PAD:7323 0.0751765
rPAD/3950 PAD:7320 PAD:13028 1.5
rPAD/3951 PAD:7319 PAD:7322 0.0751765
rPAD/3952 PAD:7319 PAD:7320 1.5
rPAD/3953 PAD:7317 PAD:13021 0.0751765
rPAD/3954 PAD:7317 PAD:7320 0.0375882
rPAD/3955 PAD:7317 PAD:13025 1.5
rPAD/3956 PAD:7316 PAD:7319 0.0375882
rPAD/3957 PAD:7316 PAD:7317 1.5
rPAD/3958 PAD:7313 PAD:7316 0.0751765
rPAD/3959 PAD:7313 PAD:13021 1.5
rPAD/3960 PAD:7311 PAD:13015 0.0751765
rPAD/3961 PAD:7311 PAD:13021 0.0375882
rPAD/3962 PAD:7311 PAD:13019 1.5
rPAD/3963 PAD:7310 PAD:7313 0.0375882
rPAD/3964 PAD:7310 PAD:7311 1.5
rPAD/3965 PAD:7307 PAD:7310 0.0751765
rPAD/3966 PAD:7307 PAD:13015 1.5
rPAD/3967 PAD:7304 PAD:7307 0.0375882
rPAD/3968 PAD:7304 PAD:13012 1.5
rPAD/3969 PAD:7301 PAD:7304 0.0751765
rPAD/3970 PAD:7301 PAD:13009 1.5
rPAD/3971 PAD:7299 PAD:13003 0.0751765
rPAD/3972 PAD:7299 PAD:13009 0.0375882
rPAD/3973 PAD:7299 PAD:13007 1.5
rPAD/3974 PAD:7298 PAD:7301 0.0375882
rPAD/3975 PAD:7298 PAD:7299 1.5
rPAD/3976 PAD:7295 PAD:7298 0.0751765
rPAD/3977 PAD:7295 PAD:13003 1.5
rPAD/3978 PAD:7292 PAD:7295 0.0375882
rPAD/3979 PAD:7292 PAD:13000 1.5
rPAD/3980 PAD:7290 PAD:13000 0.0751765
rPAD/3981 PAD:7290 PAD:12998 1.5
rPAD/3982 PAD:7289 PAD:7292 0.0751765
rPAD/3983 PAD:7289 PAD:7290 1.5
rPAD/3984 PAD:7287 PAD:7290 0.0375882
rPAD/3985 PAD:7287 PAD:12995 1.5
rPAD/3986 PAD:7286 PAD:7289 0.0375882
rPAD/3987 PAD:7286 PAD:7287 1.5
rPAD/3988 PAD:7284 PAD:7287 0.0751765
rPAD/3989 PAD:7284 PAD:12992 1.5
rPAD/3990 PAD:7283 PAD:7286 0.0751765
rPAD/3991 PAD:7283 PAD:7284 1.5
rPAD/3992 PAD:7281 PAD:7284 0.0375882
rPAD/3993 PAD:7281 PAD:12989 1.5
rPAD/3994 PAD:7280 PAD:7283 0.0375882
rPAD/3995 PAD:7280 PAD:7281 1.5
rPAD/3996 PAD:7278 PAD:7281 0.0751765
rPAD/3997 PAD:7278 PAD:12986 1.5
rPAD/3998 PAD:7277 PAD:7280 0.0751765
rPAD/3999 PAD:7277 PAD:7278 1.5
rPAD/4000 PAD:7275 PAD:12979 0.0751765
rPAD/4001 PAD:7275 PAD:7278 0.0375882
rPAD/4002 PAD:7275 PAD:12983 1.5
rPAD/4003 PAD:7274 PAD:7277 0.0375882
rPAD/4004 PAD:7274 PAD:7275 1.5
rPAD/4005 PAD:7271 PAD:7274 0.0751765
rPAD/4006 PAD:7271 PAD:12979 1.5
rPAD/4007 PAD:7269 PAD:12979 0.0375882
rPAD/4008 PAD:7269 PAD:12977 1.5
rPAD/4009 PAD:7268 PAD:7271 0.0375882
rPAD/4010 PAD:7268 PAD:7269 1.5
rPAD/4011 PAD:7266 PAD:7269 0.0751765
rPAD/4012 PAD:7266 PAD:12974 1.5
rPAD/4013 PAD:7265 PAD:7268 0.0751765
rPAD/4014 PAD:7265 PAD:7266 1.5
rPAD/4015 PAD:7263 PAD:12967 0.0751765
rPAD/4016 PAD:7263 PAD:7266 0.0375882
rPAD/4017 PAD:7263 PAD:12971 1.5
rPAD/4018 PAD:7262 PAD:7265 0.0375882
rPAD/4019 PAD:7262 PAD:7263 1.5
rPAD/4020 PAD:7259 PAD:7262 0.0751765
rPAD/4021 PAD:7259 PAD:12967 1.5
rPAD/4022 PAD:7256 PAD:7259 0.0375882
rPAD/4023 PAD:7256 PAD:12964 1.5
rPAD/4024 PAD:7253 PAD:7256 0.0751765
rPAD/4025 PAD:7253 PAD:12961 1.5
rPAD/4026 PAD:7250 PAD:7253 0.0375882
rPAD/4027 PAD:7250 PAD:12958 1.5
rPAD/4028 PAD:7247 PAD:7250 0.0751765
rPAD/4029 PAD:7247 PAD:12955 1.5
rPAD/4030 PAD:7245 PAD:12955 0.0375882
rPAD/4031 PAD:7245 PAD:12953 1.5
rPAD/4032 PAD:7244 PAD:7247 0.0375882
rPAD/4033 PAD:7244 PAD:7245 1.5
rPAD/4034 PAD:7242 PAD:12946 0.0375882
rPAD/4035 PAD:7242 PAD:7245 0.0751765
rPAD/4036 PAD:7242 PAD:12950 1.5
rPAD/4037 PAD:7241 PAD:7244 0.0751765
rPAD/4038 PAD:7241 PAD:7242 1.5
rPAD/4039 PAD:7238 PAD:7241 0.0375882
rPAD/4040 PAD:7238 PAD:12946 1.5
rPAD/4041 PAD:7236 PAD:12946 0.0751765
rPAD/4042 PAD:7236 PAD:12944 1.5
rPAD/4043 PAD:7235 PAD:7238 0.0751765
rPAD/4044 PAD:7235 PAD:7236 1.5
rPAD/4045 PAD:7233 PAD:7236 0.0375882
rPAD/4046 PAD:7233 PAD:12941 1.5
rPAD/4047 PAD:7232 PAD:7235 0.0375882
rPAD/4048 PAD:7232 PAD:7233 1.5
rPAD/4049 PAD:7230 PAD:7233 0.0751765
rPAD/4050 PAD:7230 PAD:12938 1.5
rPAD/4051 PAD:7229 PAD:7232 0.0751765
rPAD/4052 PAD:7229 PAD:7230 1.5
rPAD/4053 PAD:7227 PAD:7230 0.0375882
rPAD/4054 PAD:7227 PAD:12935 1.5
rPAD/4055 PAD:7226 PAD:7229 0.0375882
rPAD/4056 PAD:7226 PAD:7227 1.5
rPAD/4057 PAD:7224 PAD:7227 0.0751765
rPAD/4058 PAD:7224 PAD:12932 1.5
rPAD/4059 PAD:7223 PAD:7226 0.0751765
rPAD/4060 PAD:7223 PAD:7224 1.5
rPAD/4061 PAD:7221 PAD:12925 0.0751765
rPAD/4062 PAD:7221 PAD:7224 0.0375882
rPAD/4063 PAD:7221 PAD:12929 1.5
rPAD/4064 PAD:7220 PAD:7223 0.0375882
rPAD/4065 PAD:7220 PAD:7221 1.5
rPAD/4066 PAD:7217 PAD:7220 0.0751765
rPAD/4067 PAD:7217 PAD:12925 1.5
rPAD/4068 PAD:7215 PAD:12925 0.0375882
rPAD/4069 PAD:7215 PAD:12923 1.5
rPAD/4070 PAD:7214 PAD:7217 0.0375882
rPAD/4071 PAD:7214 PAD:7215 1.5
rPAD/4072 PAD:7212 PAD:7215 0.0751765
rPAD/4073 PAD:7212 PAD:12920 1.5
rPAD/4074 PAD:7211 PAD:7214 0.0751765
rPAD/4075 PAD:7211 PAD:7212 1.5
rPAD/4076 PAD:7209 PAD:7212 0.0375882
rPAD/4077 PAD:7209 PAD:12917 1.5
rPAD/4078 PAD:7208 PAD:7211 0.0375882
rPAD/4079 PAD:7208 PAD:7209 1.5
rPAD/4080 PAD:7206 PAD:7209 0.0751765
rPAD/4081 PAD:7206 PAD:12914 1.5
rPAD/4082 PAD:7205 PAD:7208 0.0751765
rPAD/4083 PAD:7205 PAD:7206 1.5
rPAD/4084 PAD:7203 PAD:7206 0.0375882
rPAD/4085 PAD:7203 PAD:12911 1.5
rPAD/4086 PAD:7202 PAD:7205 0.0375882
rPAD/4087 PAD:7202 PAD:7203 1.5
rPAD/4088 PAD:7200 PAD:7203 0.0751765
rPAD/4089 PAD:7200 PAD:12908 1.5
rPAD/4090 PAD:7199 PAD:7202 0.0751765
rPAD/4091 PAD:7199 PAD:7200 1.5
rPAD/4092 PAD:7197 PAD:7200 0.0375882
rPAD/4093 PAD:7197 PAD:12905 1.5
rPAD/4094 PAD:7196 PAD:7199 0.0375882
rPAD/4095 PAD:7196 PAD:7197 1.5
rPAD/4096 PAD:7194 PAD:14940 0.0283817
rPAD/4097 PAD:7194 PAD:7197 0.0751765
rPAD/4098 PAD:7194 PAD:12902 1.5
rPAD/4099 PAD:7193 PAD:9231 0.0378785
rPAD/4100 PAD:7193 PAD:7196 0.0751765
rPAD/4101 PAD:7193 PAD:7194 1.5
rPAD/4102 PAD:7189 PAD:12729 0.0100588
rPAD/4103 PAD:7189 PAD:12897 1.5
rPAD/4104 PAD:7188 PAD:9396 0.0670908
rPAD/4105 PAD:7188 PAD:7189 1.5
rPAD/4106 PAD:7186 PAD:7189 0.0751765
rPAD/4107 PAD:7186 PAD:12894 1.5
rPAD/4108 PAD:7185 PAD:7188 0.0751765
rPAD/4109 PAD:7185 PAD:7186 1.5
rPAD/4110 PAD:7183 PAD:12887 0.0751765
rPAD/4111 PAD:7183 PAD:7186 0.0375882
rPAD/4112 PAD:7183 PAD:12891 1.5
rPAD/4113 PAD:7182 PAD:7185 0.0375882
rPAD/4114 PAD:7182 PAD:7183 1.5
rPAD/4115 PAD:7179 PAD:7182 0.0751765
rPAD/4116 PAD:7179 PAD:12887 1.5
rPAD/4117 PAD:7177 PAD:12887 0.0375882
rPAD/4118 PAD:7177 PAD:12885 1.5
rPAD/4119 PAD:7176 PAD:7179 0.0375882
rPAD/4120 PAD:7176 PAD:7177 1.5
rPAD/4121 PAD:7174 PAD:7177 0.0751765
rPAD/4122 PAD:7174 PAD:12882 1.5
rPAD/4123 PAD:7173 PAD:7176 0.0751765
rPAD/4124 PAD:7173 PAD:7174 1.5
rPAD/4125 PAD:7171 PAD:7174 0.0375882
rPAD/4126 PAD:7171 PAD:12879 1.5
rPAD/4127 PAD:7170 PAD:7173 0.0375882
rPAD/4128 PAD:7170 PAD:7171 1.5
rPAD/4129 PAD:7168 PAD:7171 0.0751765
rPAD/4130 PAD:7168 PAD:12876 1.5
rPAD/4131 PAD:7167 PAD:7170 0.0751765
rPAD/4132 PAD:7167 PAD:7168 1.5
rPAD/4133 PAD:7165 PAD:7168 0.0375882
rPAD/4134 PAD:7165 PAD:12873 1.5
rPAD/4135 PAD:7164 PAD:7167 0.0375882
rPAD/4136 PAD:7164 PAD:7165 1.5
rPAD/4137 PAD:7162 PAD:7165 0.0751765
rPAD/4138 PAD:7162 PAD:12870 1.5
rPAD/4139 PAD:7161 PAD:7164 0.0751765
rPAD/4140 PAD:7161 PAD:7162 1.5
rPAD/4141 PAD:7159 PAD:7162 0.0375882
rPAD/4142 PAD:7159 PAD:12867 1.5
rPAD/4143 PAD:7158 PAD:7161 0.0375882
rPAD/4144 PAD:7158 PAD:7159 1.5
rPAD/4145 PAD:7156 PAD:7159 0.0751765
rPAD/4146 PAD:7156 PAD:12864 1.5
rPAD/4147 PAD:7155 PAD:7158 0.0751765
rPAD/4148 PAD:7155 PAD:7156 1.5
rPAD/4149 PAD:7153 PAD:7156 0.0375882
rPAD/4150 PAD:7153 PAD:12861 1.5
rPAD/4151 PAD:7152 PAD:7155 0.0375882
rPAD/4152 PAD:7152 PAD:7153 1.5
rPAD/4153 PAD:7150 PAD:7153 0.0751765
rPAD/4154 PAD:7150 PAD:12858 1.5
rPAD/4155 PAD:7149 PAD:7152 0.0751765
rPAD/4156 PAD:7149 PAD:7150 1.5
rPAD/4157 PAD:7147 PAD:12851 0.0751765
rPAD/4158 PAD:7147 PAD:7150 0.0375882
rPAD/4159 PAD:7147 PAD:12855 1.5
rPAD/4160 PAD:7146 PAD:7149 0.0375882
rPAD/4161 PAD:7146 PAD:7147 1.5
rPAD/4162 PAD:7143 PAD:7146 0.0751765
rPAD/4163 PAD:7143 PAD:12851 1.5
rPAD/4164 PAD:7141 PAD:12845 0.0751765
rPAD/4165 PAD:7141 PAD:12851 0.0375882
rPAD/4166 PAD:7141 PAD:12849 1.5
rPAD/4167 PAD:7140 PAD:7143 0.0375882
rPAD/4168 PAD:7140 PAD:7141 1.5
rPAD/4169 PAD:7137 PAD:7140 0.0751765
rPAD/4170 PAD:7137 PAD:12845 1.5
rPAD/4171 PAD:7134 PAD:7137 0.0375882
rPAD/4172 PAD:7134 PAD:12842 1.5
rPAD/4173 PAD:7131 PAD:7134 0.0751765
rPAD/4174 PAD:7131 PAD:12839 1.5
rPAD/4175 PAD:7129 PAD:12833 0.0751765
rPAD/4176 PAD:7129 PAD:12839 0.0375882
rPAD/4177 PAD:7129 PAD:12837 1.5
rPAD/4178 PAD:7128 PAD:7131 0.0375882
rPAD/4179 PAD:7128 PAD:7129 1.5
rPAD/4180 PAD:7125 PAD:7128 0.0751765
rPAD/4181 PAD:7125 PAD:12833 1.5
rPAD/4182 PAD:7122 PAD:7125 0.0375882
rPAD/4183 PAD:7122 PAD:12830 1.5
rPAD/4184 PAD:7120 PAD:12830 0.0751765
rPAD/4185 PAD:7120 PAD:12828 1.5
rPAD/4186 PAD:7119 PAD:7122 0.0751765
rPAD/4187 PAD:7119 PAD:7120 1.5
rPAD/4188 PAD:7117 PAD:7120 0.0375882
rPAD/4189 PAD:7117 PAD:12825 1.5
rPAD/4190 PAD:7116 PAD:7119 0.0375882
rPAD/4191 PAD:7116 PAD:7117 1.5
rPAD/4192 PAD:7114 PAD:7117 0.0751765
rPAD/4193 PAD:7114 PAD:12822 1.5
rPAD/4194 PAD:7113 PAD:7116 0.0751765
rPAD/4195 PAD:7113 PAD:7114 1.5
rPAD/4196 PAD:7111 PAD:7114 0.0375882
rPAD/4197 PAD:7111 PAD:12819 1.5
rPAD/4198 PAD:7110 PAD:7113 0.0375882
rPAD/4199 PAD:7110 PAD:7111 1.5
rPAD/4200 PAD:7108 PAD:7111 0.0751765
rPAD/4201 PAD:7108 PAD:12816 1.5
rPAD/4202 PAD:7107 PAD:7110 0.0751765
rPAD/4203 PAD:7107 PAD:7108 1.5
rPAD/4204 PAD:7105 PAD:12809 0.0751765
rPAD/4205 PAD:7105 PAD:7108 0.0375882
rPAD/4206 PAD:7105 PAD:12813 1.5
rPAD/4207 PAD:7104 PAD:7107 0.0375882
rPAD/4208 PAD:7104 PAD:7105 1.5
rPAD/4209 PAD:7101 PAD:7104 0.0751765
rPAD/4210 PAD:7101 PAD:12809 1.5
rPAD/4211 PAD:7099 PAD:12809 0.0375882
rPAD/4212 PAD:7099 PAD:12807 1.5
rPAD/4213 PAD:7098 PAD:7101 0.0375882
rPAD/4214 PAD:7098 PAD:7099 1.5
rPAD/4215 PAD:7096 PAD:7099 0.0751765
rPAD/4216 PAD:7096 PAD:12804 1.5
rPAD/4217 PAD:7095 PAD:7098 0.0751765
rPAD/4218 PAD:7095 PAD:7096 1.5
rPAD/4219 PAD:7093 PAD:12797 0.0751765
rPAD/4220 PAD:7093 PAD:7096 0.0375882
rPAD/4221 PAD:7093 PAD:12801 1.5
rPAD/4222 PAD:7092 PAD:7095 0.0375882
rPAD/4223 PAD:7092 PAD:7093 1.5
rPAD/4224 PAD:7089 PAD:7092 0.0751765
rPAD/4225 PAD:7089 PAD:12797 1.5
rPAD/4226 PAD:7086 PAD:7089 0.0375882
rPAD/4227 PAD:7086 PAD:12794 1.5
rPAD/4228 PAD:7083 PAD:7086 0.0751765
rPAD/4229 PAD:7083 PAD:12791 1.5
rPAD/4230 PAD:7080 PAD:7083 0.0375882
rPAD/4231 PAD:7080 PAD:12788 1.5
rPAD/4232 PAD:7077 PAD:7080 0.0751765
rPAD/4233 PAD:7077 PAD:12785 1.5
rPAD/4234 PAD:7075 PAD:12785 0.0375882
rPAD/4235 PAD:7075 PAD:12783 1.5
rPAD/4236 PAD:7074 PAD:7077 0.0375882
rPAD/4237 PAD:7074 PAD:7075 1.5
rPAD/4238 PAD:7072 PAD:12776 0.0375882
rPAD/4239 PAD:7072 PAD:7075 0.0751765
rPAD/4240 PAD:7072 PAD:12780 1.5
rPAD/4241 PAD:7071 PAD:7074 0.0751765
rPAD/4242 PAD:7071 PAD:7072 1.5
rPAD/4243 PAD:7068 PAD:7071 0.0375882
rPAD/4244 PAD:7068 PAD:12776 1.5
rPAD/4245 PAD:7066 PAD:12776 0.0751765
rPAD/4246 PAD:7066 PAD:12774 1.5
rPAD/4247 PAD:7065 PAD:7068 0.0751765
rPAD/4248 PAD:7065 PAD:7066 1.5
rPAD/4249 PAD:7063 PAD:7066 0.0375882
rPAD/4250 PAD:7063 PAD:12771 1.5
rPAD/4251 PAD:7062 PAD:7065 0.0375882
rPAD/4252 PAD:7062 PAD:7063 1.5
rPAD/4253 PAD:7060 PAD:7063 0.0751765
rPAD/4254 PAD:7060 PAD:12768 1.5
rPAD/4255 PAD:7059 PAD:7062 0.0751765
rPAD/4256 PAD:7059 PAD:7060 1.5
rPAD/4257 PAD:7057 PAD:7060 0.0375882
rPAD/4258 PAD:7057 PAD:12765 1.5
rPAD/4259 PAD:7056 PAD:7059 0.0375882
rPAD/4260 PAD:7056 PAD:7057 1.5
rPAD/4261 PAD:7054 PAD:7057 0.0751765
rPAD/4262 PAD:7054 PAD:12762 1.5
rPAD/4263 PAD:7053 PAD:7056 0.0751765
rPAD/4264 PAD:7053 PAD:7054 1.5
rPAD/4265 PAD:7051 PAD:12755 0.0751765
rPAD/4266 PAD:7051 PAD:7054 0.0375882
rPAD/4267 PAD:7051 PAD:12759 1.5
rPAD/4268 PAD:7050 PAD:7053 0.0375882
rPAD/4269 PAD:7050 PAD:7051 1.5
rPAD/4270 PAD:7047 PAD:7050 0.0751765
rPAD/4271 PAD:7047 PAD:12755 1.5
rPAD/4272 PAD:7045 PAD:12755 0.0375882
rPAD/4273 PAD:7045 PAD:12753 1.5
rPAD/4274 PAD:7044 PAD:7047 0.0375882
rPAD/4275 PAD:7044 PAD:7045 1.5
rPAD/4276 PAD:7042 PAD:7045 0.0751765
rPAD/4277 PAD:7042 PAD:12750 1.5
rPAD/4278 PAD:7041 PAD:7044 0.0751765
rPAD/4279 PAD:7041 PAD:7042 1.5
rPAD/4280 PAD:7039 PAD:7042 0.0375882
rPAD/4281 PAD:7039 PAD:12747 1.5
rPAD/4282 PAD:7038 PAD:7041 0.0375882
rPAD/4283 PAD:7038 PAD:7039 1.5
rPAD/4284 PAD:7036 PAD:7039 0.0751765
rPAD/4285 PAD:7036 PAD:12744 1.5
rPAD/4286 PAD:7035 PAD:7038 0.0751765
rPAD/4287 PAD:7035 PAD:7036 1.5
rPAD/4288 PAD:7033 PAD:7036 0.0375882
rPAD/4289 PAD:7033 PAD:12741 1.5
rPAD/4290 PAD:7032 PAD:7035 0.0375882
rPAD/4291 PAD:7032 PAD:7033 1.5
rPAD/4292 PAD:7030 PAD:7033 0.0751765
rPAD/4293 PAD:7030 PAD:12738 1.5
rPAD/4294 PAD:7029 PAD:7032 0.0751765
rPAD/4295 PAD:7029 PAD:7030 1.5
rPAD/4296 PAD:7027 PAD:7030 0.0375882
rPAD/4297 PAD:7027 PAD:12735 1.5
rPAD/4298 PAD:7026 PAD:7029 0.0375882
rPAD/4299 PAD:7026 PAD:7027 1.5
rPAD/4300 PAD:7024 PAD:14935 0.0283817
rPAD/4301 PAD:7024 PAD:7027 0.0751765
rPAD/4302 PAD:7024 PAD:12732 1.5
rPAD/4303 PAD:7023 PAD:9224 0.0378785
rPAD/4304 PAD:7023 PAD:7026 0.0751765
rPAD/4305 PAD:7023 PAD:7024 1.5
rPAD/4306 PAD:7019 PAD:12559 0.0100588
rPAD/4307 PAD:7019 PAD:12727 1.5
rPAD/4308 PAD:7018 PAD:9392 0.0670908
rPAD/4309 PAD:7018 PAD:7019 1.5
rPAD/4310 PAD:7016 PAD:7019 0.0751765
rPAD/4311 PAD:7016 PAD:12724 1.5
rPAD/4312 PAD:7015 PAD:7018 0.0751765
rPAD/4313 PAD:7015 PAD:7016 1.5
rPAD/4314 PAD:7013 PAD:12717 0.0751765
rPAD/4315 PAD:7013 PAD:7016 0.0375882
rPAD/4316 PAD:7013 PAD:12721 1.5
rPAD/4317 PAD:7012 PAD:7015 0.0375882
rPAD/4318 PAD:7012 PAD:7013 1.5
rPAD/4319 PAD:7009 PAD:7012 0.0751765
rPAD/4320 PAD:7009 PAD:12717 1.5
rPAD/4321 PAD:7007 PAD:12717 0.0375882
rPAD/4322 PAD:7007 PAD:12715 1.5
rPAD/4323 PAD:7006 PAD:7009 0.0375882
rPAD/4324 PAD:7006 PAD:7007 1.5
rPAD/4325 PAD:7004 PAD:7007 0.0751765
rPAD/4326 PAD:7004 PAD:12712 1.5
rPAD/4327 PAD:7003 PAD:7006 0.0751765
rPAD/4328 PAD:7003 PAD:7004 1.5
rPAD/4329 PAD:7001 PAD:7004 0.0375882
rPAD/4330 PAD:7001 PAD:12709 1.5
rPAD/4331 PAD:7000 PAD:7003 0.0375882
rPAD/4332 PAD:7000 PAD:7001 1.5
rPAD/4333 PAD:6998 PAD:7001 0.0751765
rPAD/4334 PAD:6998 PAD:12706 1.5
rPAD/4335 PAD:6997 PAD:7000 0.0751765
rPAD/4336 PAD:6997 PAD:6998 1.5
rPAD/4337 PAD:6995 PAD:6998 0.0375882
rPAD/4338 PAD:6995 PAD:12703 1.5
rPAD/4339 PAD:6994 PAD:6997 0.0375882
rPAD/4340 PAD:6994 PAD:6995 1.5
rPAD/4341 PAD:6992 PAD:6995 0.0751765
rPAD/4342 PAD:6992 PAD:12700 1.5
rPAD/4343 PAD:6991 PAD:6994 0.0751765
rPAD/4344 PAD:6991 PAD:6992 1.5
rPAD/4345 PAD:6989 PAD:6992 0.0375882
rPAD/4346 PAD:6989 PAD:12697 1.5
rPAD/4347 PAD:6988 PAD:6991 0.0375882
rPAD/4348 PAD:6988 PAD:6989 1.5
rPAD/4349 PAD:6986 PAD:6989 0.0751765
rPAD/4350 PAD:6986 PAD:12694 1.5
rPAD/4351 PAD:6985 PAD:6988 0.0751765
rPAD/4352 PAD:6985 PAD:6986 1.5
rPAD/4353 PAD:6983 PAD:6986 0.0375882
rPAD/4354 PAD:6983 PAD:12691 1.5
rPAD/4355 PAD:6982 PAD:6985 0.0375882
rPAD/4356 PAD:6982 PAD:6983 1.5
rPAD/4357 PAD:6980 PAD:6983 0.0751765
rPAD/4358 PAD:6980 PAD:12688 1.5
rPAD/4359 PAD:6979 PAD:6982 0.0751765
rPAD/4360 PAD:6979 PAD:6980 1.5
rPAD/4361 PAD:6977 PAD:12681 0.0751765
rPAD/4362 PAD:6977 PAD:6980 0.0375882
rPAD/4363 PAD:6977 PAD:12685 1.5
rPAD/4364 PAD:6976 PAD:6979 0.0375882
rPAD/4365 PAD:6976 PAD:6977 1.5
rPAD/4366 PAD:6973 PAD:6976 0.0751765
rPAD/4367 PAD:6973 PAD:12681 1.5
rPAD/4368 PAD:6971 PAD:12675 0.0751765
rPAD/4369 PAD:6971 PAD:12681 0.0375882
rPAD/4370 PAD:6971 PAD:12679 1.5
rPAD/4371 PAD:6970 PAD:6973 0.0375882
rPAD/4372 PAD:6970 PAD:6971 1.5
rPAD/4373 PAD:6967 PAD:6970 0.0751765
rPAD/4374 PAD:6967 PAD:12675 1.5
rPAD/4375 PAD:6964 PAD:6967 0.0375882
rPAD/4376 PAD:6964 PAD:12672 1.5
rPAD/4377 PAD:6961 PAD:6964 0.0751765
rPAD/4378 PAD:6961 PAD:12669 1.5
rPAD/4379 PAD:6959 PAD:12663 0.0751765
rPAD/4380 PAD:6959 PAD:12669 0.0375882
rPAD/4381 PAD:6959 PAD:12667 1.5
rPAD/4382 PAD:6958 PAD:6961 0.0375882
rPAD/4383 PAD:6958 PAD:6959 1.5
rPAD/4384 PAD:6955 PAD:6958 0.0751765
rPAD/4385 PAD:6955 PAD:12663 1.5
rPAD/4386 PAD:6952 PAD:6955 0.0375882
rPAD/4387 PAD:6952 PAD:12660 1.5
rPAD/4388 PAD:6950 PAD:12660 0.0751765
rPAD/4389 PAD:6950 PAD:12658 1.5
rPAD/4390 PAD:6949 PAD:6952 0.0751765
rPAD/4391 PAD:6949 PAD:6950 1.5
rPAD/4392 PAD:6947 PAD:6950 0.0375882
rPAD/4393 PAD:6947 PAD:12655 1.5
rPAD/4394 PAD:6946 PAD:6949 0.0375882
rPAD/4395 PAD:6946 PAD:6947 1.5
rPAD/4396 PAD:6944 PAD:6947 0.0751765
rPAD/4397 PAD:6944 PAD:12652 1.5
rPAD/4398 PAD:6943 PAD:6946 0.0751765
rPAD/4399 PAD:6943 PAD:6944 1.5
rPAD/4400 PAD:6941 PAD:6944 0.0375882
rPAD/4401 PAD:6941 PAD:12649 1.5
rPAD/4402 PAD:6940 PAD:6943 0.0375882
rPAD/4403 PAD:6940 PAD:6941 1.5
rPAD/4404 PAD:6938 PAD:6941 0.0751765
rPAD/4405 PAD:6938 PAD:12646 1.5
rPAD/4406 PAD:6937 PAD:6940 0.0751765
rPAD/4407 PAD:6937 PAD:6938 1.5
rPAD/4408 PAD:6935 PAD:12639 0.0751765
rPAD/4409 PAD:6935 PAD:6938 0.0375882
rPAD/4410 PAD:6935 PAD:12643 1.5
rPAD/4411 PAD:6934 PAD:6937 0.0375882
rPAD/4412 PAD:6934 PAD:6935 1.5
rPAD/4413 PAD:6931 PAD:6934 0.0751765
rPAD/4414 PAD:6931 PAD:12639 1.5
rPAD/4415 PAD:6929 PAD:12639 0.0375882
rPAD/4416 PAD:6929 PAD:12637 1.5
rPAD/4417 PAD:6928 PAD:6931 0.0375882
rPAD/4418 PAD:6928 PAD:6929 1.5
rPAD/4419 PAD:6926 PAD:6929 0.0751765
rPAD/4420 PAD:6926 PAD:12634 1.5
rPAD/4421 PAD:6925 PAD:6928 0.0751765
rPAD/4422 PAD:6925 PAD:6926 1.5
rPAD/4423 PAD:6923 PAD:12627 0.0751765
rPAD/4424 PAD:6923 PAD:6926 0.0375882
rPAD/4425 PAD:6923 PAD:12631 1.5
rPAD/4426 PAD:6922 PAD:6925 0.0375882
rPAD/4427 PAD:6922 PAD:6923 1.5
rPAD/4428 PAD:6919 PAD:6922 0.0751765
rPAD/4429 PAD:6919 PAD:12627 1.5
rPAD/4430 PAD:6916 PAD:6919 0.0375882
rPAD/4431 PAD:6916 PAD:12624 1.5
rPAD/4432 PAD:6913 PAD:6916 0.0751765
rPAD/4433 PAD:6913 PAD:12621 1.5
rPAD/4434 PAD:6910 PAD:6913 0.0375882
rPAD/4435 PAD:6910 PAD:12618 1.5
rPAD/4436 PAD:6907 PAD:6910 0.0751765
rPAD/4437 PAD:6907 PAD:12615 1.5
rPAD/4438 PAD:6905 PAD:12615 0.0375882
rPAD/4439 PAD:6905 PAD:12613 1.5
rPAD/4440 PAD:6904 PAD:6907 0.0375882
rPAD/4441 PAD:6904 PAD:6905 1.5
rPAD/4442 PAD:6902 PAD:12606 0.0375882
rPAD/4443 PAD:6902 PAD:6905 0.0751765
rPAD/4444 PAD:6902 PAD:12610 1.5
rPAD/4445 PAD:6901 PAD:6904 0.0751765
rPAD/4446 PAD:6901 PAD:6902 1.5
rPAD/4447 PAD:6898 PAD:6901 0.0375882
rPAD/4448 PAD:6898 PAD:12606 1.5
rPAD/4449 PAD:6896 PAD:12606 0.0751765
rPAD/4450 PAD:6896 PAD:12604 1.5
rPAD/4451 PAD:6895 PAD:6898 0.0751765
rPAD/4452 PAD:6895 PAD:6896 1.5
rPAD/4453 PAD:6893 PAD:6896 0.0375882
rPAD/4454 PAD:6893 PAD:12601 1.5
rPAD/4455 PAD:6892 PAD:6895 0.0375882
rPAD/4456 PAD:6892 PAD:6893 1.5
rPAD/4457 PAD:6890 PAD:6893 0.0751765
rPAD/4458 PAD:6890 PAD:12598 1.5
rPAD/4459 PAD:6889 PAD:6892 0.0751765
rPAD/4460 PAD:6889 PAD:6890 1.5
rPAD/4461 PAD:6887 PAD:6890 0.0375882
rPAD/4462 PAD:6887 PAD:12595 1.5
rPAD/4463 PAD:6886 PAD:6889 0.0375882
rPAD/4464 PAD:6886 PAD:6887 1.5
rPAD/4465 PAD:6884 PAD:6887 0.0751765
rPAD/4466 PAD:6884 PAD:12592 1.5
rPAD/4467 PAD:6883 PAD:6886 0.0751765
rPAD/4468 PAD:6883 PAD:6884 1.5
rPAD/4469 PAD:6881 PAD:12585 0.0751765
rPAD/4470 PAD:6881 PAD:6884 0.0375882
rPAD/4471 PAD:6881 PAD:12589 1.5
rPAD/4472 PAD:6880 PAD:6883 0.0375882
rPAD/4473 PAD:6880 PAD:6881 1.5
rPAD/4474 PAD:6877 PAD:6880 0.0751765
rPAD/4475 PAD:6877 PAD:12585 1.5
rPAD/4476 PAD:6875 PAD:12585 0.0375882
rPAD/4477 PAD:6875 PAD:12583 1.5
rPAD/4478 PAD:6874 PAD:6877 0.0375882
rPAD/4479 PAD:6874 PAD:6875 1.5
rPAD/4480 PAD:6872 PAD:6875 0.0751765
rPAD/4481 PAD:6872 PAD:12580 1.5
rPAD/4482 PAD:6871 PAD:6874 0.0751765
rPAD/4483 PAD:6871 PAD:6872 1.5
rPAD/4484 PAD:6869 PAD:6872 0.0375882
rPAD/4485 PAD:6869 PAD:12577 1.5
rPAD/4486 PAD:6868 PAD:6871 0.0375882
rPAD/4487 PAD:6868 PAD:6869 1.5
rPAD/4488 PAD:6866 PAD:6869 0.0751765
rPAD/4489 PAD:6866 PAD:12574 1.5
rPAD/4490 PAD:6865 PAD:6868 0.0751765
rPAD/4491 PAD:6865 PAD:6866 1.5
rPAD/4492 PAD:6863 PAD:6866 0.0375882
rPAD/4493 PAD:6863 PAD:12571 1.5
rPAD/4494 PAD:6862 PAD:6865 0.0375882
rPAD/4495 PAD:6862 PAD:6863 1.5
rPAD/4496 PAD:6860 PAD:6863 0.0751765
rPAD/4497 PAD:6860 PAD:12568 1.5
rPAD/4498 PAD:6859 PAD:6862 0.0751765
rPAD/4499 PAD:6859 PAD:6860 1.5
rPAD/4500 PAD:6857 PAD:6860 0.0375882
rPAD/4501 PAD:6857 PAD:12565 1.5
rPAD/4502 PAD:6856 PAD:6859 0.0375882
rPAD/4503 PAD:6856 PAD:6857 1.5
rPAD/4504 PAD:6854 PAD:14927 0.0283817
rPAD/4505 PAD:6854 PAD:6857 0.0751765
rPAD/4506 PAD:6854 PAD:12562 1.5
rPAD/4507 PAD:6853 PAD:9217 0.0378785
rPAD/4508 PAD:6853 PAD:6856 0.0751765
rPAD/4509 PAD:6853 PAD:6854 1.5
rPAD/4510 PAD:6849 PAD:12389 0.0100588
rPAD/4511 PAD:6849 PAD:12557 1.5
rPAD/4512 PAD:6848 PAD:9388 0.0670908
rPAD/4513 PAD:6848 PAD:6849 1.5
rPAD/4514 PAD:6846 PAD:6849 0.0751765
rPAD/4515 PAD:6846 PAD:12554 1.5
rPAD/4516 PAD:6845 PAD:6848 0.0751765
rPAD/4517 PAD:6845 PAD:6846 1.5
rPAD/4518 PAD:6843 PAD:12547 0.0751765
rPAD/4519 PAD:6843 PAD:6846 0.0375882
rPAD/4520 PAD:6843 PAD:12551 1.5
rPAD/4521 PAD:6842 PAD:6845 0.0375882
rPAD/4522 PAD:6842 PAD:6843 1.5
rPAD/4523 PAD:6839 PAD:6842 0.0751765
rPAD/4524 PAD:6839 PAD:12547 1.5
rPAD/4525 PAD:6837 PAD:12547 0.0375882
rPAD/4526 PAD:6837 PAD:12545 1.5
rPAD/4527 PAD:6836 PAD:6839 0.0375882
rPAD/4528 PAD:6836 PAD:6837 1.5
rPAD/4529 PAD:6834 PAD:6837 0.0751765
rPAD/4530 PAD:6834 PAD:12542 1.5
rPAD/4531 PAD:6833 PAD:6836 0.0751765
rPAD/4532 PAD:6833 PAD:6834 1.5
rPAD/4533 PAD:6831 PAD:6834 0.0375882
rPAD/4534 PAD:6831 PAD:12539 1.5
rPAD/4535 PAD:6830 PAD:6833 0.0375882
rPAD/4536 PAD:6830 PAD:6831 1.5
rPAD/4537 PAD:6828 PAD:6831 0.0751765
rPAD/4538 PAD:6828 PAD:12536 1.5
rPAD/4539 PAD:6827 PAD:6830 0.0751765
rPAD/4540 PAD:6827 PAD:6828 1.5
rPAD/4541 PAD:6825 PAD:6828 0.0375882
rPAD/4542 PAD:6825 PAD:12533 1.5
rPAD/4543 PAD:6824 PAD:6827 0.0375882
rPAD/4544 PAD:6824 PAD:6825 1.5
rPAD/4545 PAD:6822 PAD:6825 0.0751765
rPAD/4546 PAD:6822 PAD:12530 1.5
rPAD/4547 PAD:6821 PAD:6824 0.0751765
rPAD/4548 PAD:6821 PAD:6822 1.5
rPAD/4549 PAD:6819 PAD:6822 0.0375882
rPAD/4550 PAD:6819 PAD:12527 1.5
rPAD/4551 PAD:6818 PAD:6821 0.0375882
rPAD/4552 PAD:6818 PAD:6819 1.5
rPAD/4553 PAD:6816 PAD:6819 0.0751765
rPAD/4554 PAD:6816 PAD:12524 1.5
rPAD/4555 PAD:6815 PAD:6818 0.0751765
rPAD/4556 PAD:6815 PAD:6816 1.5
rPAD/4557 PAD:6813 PAD:6816 0.0375882
rPAD/4558 PAD:6813 PAD:12521 1.5
rPAD/4559 PAD:6812 PAD:6815 0.0375882
rPAD/4560 PAD:6812 PAD:6813 1.5
rPAD/4561 PAD:6810 PAD:6813 0.0751765
rPAD/4562 PAD:6810 PAD:12518 1.5
rPAD/4563 PAD:6809 PAD:6812 0.0751765
rPAD/4564 PAD:6809 PAD:6810 1.5
rPAD/4565 PAD:6807 PAD:12511 0.0751765
rPAD/4566 PAD:6807 PAD:6810 0.0375882
rPAD/4567 PAD:6807 PAD:12515 1.5
rPAD/4568 PAD:6806 PAD:6809 0.0375882
rPAD/4569 PAD:6806 PAD:6807 1.5
rPAD/4570 PAD:6803 PAD:6806 0.0751765
rPAD/4571 PAD:6803 PAD:12511 1.5
rPAD/4572 PAD:6801 PAD:12505 0.0751765
rPAD/4573 PAD:6801 PAD:12511 0.0375882
rPAD/4574 PAD:6801 PAD:12509 1.5
rPAD/4575 PAD:6800 PAD:6803 0.0375882
rPAD/4576 PAD:6800 PAD:6801 1.5
rPAD/4577 PAD:6797 PAD:6800 0.0751765
rPAD/4578 PAD:6797 PAD:12505 1.5
rPAD/4579 PAD:6794 PAD:6797 0.0375882
rPAD/4580 PAD:6794 PAD:12502 1.5
rPAD/4581 PAD:6791 PAD:6794 0.0751765
rPAD/4582 PAD:6791 PAD:12499 1.5
rPAD/4583 PAD:6789 PAD:12493 0.0751765
rPAD/4584 PAD:6789 PAD:12499 0.0375882
rPAD/4585 PAD:6789 PAD:12497 1.5
rPAD/4586 PAD:6788 PAD:6791 0.0375882
rPAD/4587 PAD:6788 PAD:6789 1.5
rPAD/4588 PAD:6785 PAD:6788 0.0751765
rPAD/4589 PAD:6785 PAD:12493 1.5
rPAD/4590 PAD:6782 PAD:6785 0.0375882
rPAD/4591 PAD:6782 PAD:12490 1.5
rPAD/4592 PAD:6780 PAD:12490 0.0751765
rPAD/4593 PAD:6780 PAD:12488 1.5
rPAD/4594 PAD:6779 PAD:6782 0.0751765
rPAD/4595 PAD:6779 PAD:6780 1.5
rPAD/4596 PAD:6777 PAD:6780 0.0375882
rPAD/4597 PAD:6777 PAD:12485 1.5
rPAD/4598 PAD:6776 PAD:6779 0.0375882
rPAD/4599 PAD:6776 PAD:6777 1.5
rPAD/4600 PAD:6774 PAD:6777 0.0751765
rPAD/4601 PAD:6774 PAD:12482 1.5
rPAD/4602 PAD:6773 PAD:6776 0.0751765
rPAD/4603 PAD:6773 PAD:6774 1.5
rPAD/4604 PAD:6771 PAD:6774 0.0375882
rPAD/4605 PAD:6771 PAD:12479 1.5
rPAD/4606 PAD:6770 PAD:6773 0.0375882
rPAD/4607 PAD:6770 PAD:6771 1.5
rPAD/4608 PAD:6768 PAD:6771 0.0751765
rPAD/4609 PAD:6768 PAD:12476 1.5
rPAD/4610 PAD:6767 PAD:6770 0.0751765
rPAD/4611 PAD:6767 PAD:6768 1.5
rPAD/4612 PAD:6765 PAD:12469 0.0751765
rPAD/4613 PAD:6765 PAD:6768 0.0375882
rPAD/4614 PAD:6765 PAD:12473 1.5
rPAD/4615 PAD:6764 PAD:6767 0.0375882
rPAD/4616 PAD:6764 PAD:6765 1.5
rPAD/4617 PAD:6761 PAD:6764 0.0751765
rPAD/4618 PAD:6761 PAD:12469 1.5
rPAD/4619 PAD:6759 PAD:12469 0.0375882
rPAD/4620 PAD:6759 PAD:12467 1.5
rPAD/4621 PAD:6758 PAD:6761 0.0375882
rPAD/4622 PAD:6758 PAD:6759 1.5
rPAD/4623 PAD:6756 PAD:6759 0.0751765
rPAD/4624 PAD:6756 PAD:12464 1.5
rPAD/4625 PAD:6755 PAD:6758 0.0751765
rPAD/4626 PAD:6755 PAD:6756 1.5
rPAD/4627 PAD:6753 PAD:12457 0.0751765
rPAD/4628 PAD:6753 PAD:6756 0.0375882
rPAD/4629 PAD:6753 PAD:12461 1.5
rPAD/4630 PAD:6752 PAD:6755 0.0375882
rPAD/4631 PAD:6752 PAD:6753 1.5
rPAD/4632 PAD:6749 PAD:6752 0.0751765
rPAD/4633 PAD:6749 PAD:12457 1.5
rPAD/4634 PAD:6746 PAD:6749 0.0375882
rPAD/4635 PAD:6746 PAD:12454 1.5
rPAD/4636 PAD:6743 PAD:6746 0.0751765
rPAD/4637 PAD:6743 PAD:12451 1.5
rPAD/4638 PAD:6740 PAD:6743 0.0375882
rPAD/4639 PAD:6740 PAD:12448 1.5
rPAD/4640 PAD:6737 PAD:6740 0.0751765
rPAD/4641 PAD:6737 PAD:12445 1.5
rPAD/4642 PAD:6735 PAD:12445 0.0375882
rPAD/4643 PAD:6735 PAD:12443 1.5
rPAD/4644 PAD:6734 PAD:6737 0.0375882
rPAD/4645 PAD:6734 PAD:6735 1.5
rPAD/4646 PAD:6732 PAD:12436 0.0375882
rPAD/4647 PAD:6732 PAD:6735 0.0751765
rPAD/4648 PAD:6732 PAD:12440 1.5
rPAD/4649 PAD:6731 PAD:6734 0.0751765
rPAD/4650 PAD:6731 PAD:6732 1.5
rPAD/4651 PAD:6728 PAD:6731 0.0375882
rPAD/4652 PAD:6728 PAD:12436 1.5
rPAD/4653 PAD:6726 PAD:12436 0.0751765
rPAD/4654 PAD:6726 PAD:12434 1.5
rPAD/4655 PAD:6725 PAD:6728 0.0751765
rPAD/4656 PAD:6725 PAD:6726 1.5
rPAD/4657 PAD:6723 PAD:6726 0.0375882
rPAD/4658 PAD:6723 PAD:12431 1.5
rPAD/4659 PAD:6722 PAD:6725 0.0375882
rPAD/4660 PAD:6722 PAD:6723 1.5
rPAD/4661 PAD:6720 PAD:6723 0.0751765
rPAD/4662 PAD:6720 PAD:12428 1.5
rPAD/4663 PAD:6719 PAD:6722 0.0751765
rPAD/4664 PAD:6719 PAD:6720 1.5
rPAD/4665 PAD:6717 PAD:6720 0.0375882
rPAD/4666 PAD:6717 PAD:12425 1.5
rPAD/4667 PAD:6716 PAD:6719 0.0375882
rPAD/4668 PAD:6716 PAD:6717 1.5
rPAD/4669 PAD:6714 PAD:6717 0.0751765
rPAD/4670 PAD:6714 PAD:12422 1.5
rPAD/4671 PAD:6713 PAD:6716 0.0751765
rPAD/4672 PAD:6713 PAD:6714 1.5
rPAD/4673 PAD:6711 PAD:12415 0.0751765
rPAD/4674 PAD:6711 PAD:6714 0.0375882
rPAD/4675 PAD:6711 PAD:12419 1.5
rPAD/4676 PAD:6710 PAD:6713 0.0375882
rPAD/4677 PAD:6710 PAD:6711 1.5
rPAD/4678 PAD:6707 PAD:6710 0.0751765
rPAD/4679 PAD:6707 PAD:12415 1.5
rPAD/4680 PAD:6705 PAD:12415 0.0375882
rPAD/4681 PAD:6705 PAD:12413 1.5
rPAD/4682 PAD:6704 PAD:6707 0.0375882
rPAD/4683 PAD:6704 PAD:6705 1.5
rPAD/4684 PAD:6702 PAD:6705 0.0751765
rPAD/4685 PAD:6702 PAD:12410 1.5
rPAD/4686 PAD:6701 PAD:6704 0.0751765
rPAD/4687 PAD:6701 PAD:6702 1.5
rPAD/4688 PAD:6699 PAD:6702 0.0375882
rPAD/4689 PAD:6699 PAD:12407 1.5
rPAD/4690 PAD:6698 PAD:6701 0.0375882
rPAD/4691 PAD:6698 PAD:6699 1.5
rPAD/4692 PAD:6696 PAD:6699 0.0751765
rPAD/4693 PAD:6696 PAD:12404 1.5
rPAD/4694 PAD:6695 PAD:6698 0.0751765
rPAD/4695 PAD:6695 PAD:6696 1.5
rPAD/4696 PAD:6693 PAD:6696 0.0375882
rPAD/4697 PAD:6693 PAD:12401 1.5
rPAD/4698 PAD:6692 PAD:6695 0.0375882
rPAD/4699 PAD:6692 PAD:6693 1.5
rPAD/4700 PAD:6690 PAD:6693 0.0751765
rPAD/4701 PAD:6690 PAD:12398 1.5
rPAD/4702 PAD:6689 PAD:6692 0.0751765
rPAD/4703 PAD:6689 PAD:6690 1.5
rPAD/4704 PAD:6687 PAD:6690 0.0375882
rPAD/4705 PAD:6687 PAD:12395 1.5
rPAD/4706 PAD:6686 PAD:6689 0.0375882
rPAD/4707 PAD:6686 PAD:6687 1.5
rPAD/4708 PAD:6684 PAD:14921 0.0283817
rPAD/4709 PAD:6684 PAD:6687 0.0751765
rPAD/4710 PAD:6684 PAD:12392 1.5
rPAD/4711 PAD:6683 PAD:9210 0.0378785
rPAD/4712 PAD:6683 PAD:6686 0.0751765
rPAD/4713 PAD:6683 PAD:6684 1.5
rPAD/4714 PAD:6679 PAD:12219 0.0100588
rPAD/4715 PAD:6679 PAD:12387 1.5
rPAD/4716 PAD:6678 PAD:9383 0.0670908
rPAD/4717 PAD:6678 PAD:6679 1.5
rPAD/4718 PAD:6676 PAD:6679 0.0751765
rPAD/4719 PAD:6676 PAD:12384 1.5
rPAD/4720 PAD:6675 PAD:6678 0.0751765
rPAD/4721 PAD:6675 PAD:6676 1.5
rPAD/4722 PAD:6673 PAD:12377 0.0751765
rPAD/4723 PAD:6673 PAD:6676 0.0375882
rPAD/4724 PAD:6673 PAD:12381 1.5
rPAD/4725 PAD:6672 PAD:6675 0.0375882
rPAD/4726 PAD:6672 PAD:6673 1.5
rPAD/4727 PAD:6669 PAD:6672 0.0751765
rPAD/4728 PAD:6669 PAD:12377 1.5
rPAD/4729 PAD:6667 PAD:12377 0.0375882
rPAD/4730 PAD:6667 PAD:12375 1.5
rPAD/4731 PAD:6666 PAD:6669 0.0375882
rPAD/4732 PAD:6666 PAD:6667 1.5
rPAD/4733 PAD:6664 PAD:6667 0.0751765
rPAD/4734 PAD:6664 PAD:12372 1.5
rPAD/4735 PAD:6663 PAD:6666 0.0751765
rPAD/4736 PAD:6663 PAD:6664 1.5
rPAD/4737 PAD:6661 PAD:6664 0.0375882
rPAD/4738 PAD:6661 PAD:12369 1.5
rPAD/4739 PAD:6660 PAD:6663 0.0375882
rPAD/4740 PAD:6660 PAD:6661 1.5
rPAD/4741 PAD:6658 PAD:6661 0.0751765
rPAD/4742 PAD:6658 PAD:12366 1.5
rPAD/4743 PAD:6657 PAD:6660 0.0751765
rPAD/4744 PAD:6657 PAD:6658 1.5
rPAD/4745 PAD:6655 PAD:6658 0.0375882
rPAD/4746 PAD:6655 PAD:12363 1.5
rPAD/4747 PAD:6654 PAD:6657 0.0375882
rPAD/4748 PAD:6654 PAD:6655 1.5
rPAD/4749 PAD:6652 PAD:6655 0.0751765
rPAD/4750 PAD:6652 PAD:12360 1.5
rPAD/4751 PAD:6651 PAD:6654 0.0751765
rPAD/4752 PAD:6651 PAD:6652 1.5
rPAD/4753 PAD:6649 PAD:6652 0.0375882
rPAD/4754 PAD:6649 PAD:12357 1.5
rPAD/4755 PAD:6648 PAD:6651 0.0375882
rPAD/4756 PAD:6648 PAD:6649 1.5
rPAD/4757 PAD:6646 PAD:6649 0.0751765
rPAD/4758 PAD:6646 PAD:12354 1.5
rPAD/4759 PAD:6645 PAD:6648 0.0751765
rPAD/4760 PAD:6645 PAD:6646 1.5
rPAD/4761 PAD:6643 PAD:6646 0.0375882
rPAD/4762 PAD:6643 PAD:12351 1.5
rPAD/4763 PAD:6642 PAD:6645 0.0375882
rPAD/4764 PAD:6642 PAD:6643 1.5
rPAD/4765 PAD:6640 PAD:6643 0.0751765
rPAD/4766 PAD:6640 PAD:12348 1.5
rPAD/4767 PAD:6639 PAD:6642 0.0751765
rPAD/4768 PAD:6639 PAD:6640 1.5
rPAD/4769 PAD:6637 PAD:12341 0.0751765
rPAD/4770 PAD:6637 PAD:6640 0.0375882
rPAD/4771 PAD:6637 PAD:12345 1.5
rPAD/4772 PAD:6636 PAD:6639 0.0375882
rPAD/4773 PAD:6636 PAD:6637 1.5
rPAD/4774 PAD:6633 PAD:6636 0.0751765
rPAD/4775 PAD:6633 PAD:12341 1.5
rPAD/4776 PAD:6631 PAD:12335 0.0751765
rPAD/4777 PAD:6631 PAD:12341 0.0375882
rPAD/4778 PAD:6631 PAD:12339 1.5
rPAD/4779 PAD:6630 PAD:6633 0.0375882
rPAD/4780 PAD:6630 PAD:6631 1.5
rPAD/4781 PAD:6627 PAD:6630 0.0751765
rPAD/4782 PAD:6627 PAD:12335 1.5
rPAD/4783 PAD:6624 PAD:6627 0.0375882
rPAD/4784 PAD:6624 PAD:12332 1.5
rPAD/4785 PAD:6621 PAD:6624 0.0751765
rPAD/4786 PAD:6621 PAD:12329 1.5
rPAD/4787 PAD:6619 PAD:12323 0.0751765
rPAD/4788 PAD:6619 PAD:12329 0.0375882
rPAD/4789 PAD:6619 PAD:12327 1.5
rPAD/4790 PAD:6618 PAD:6621 0.0375882
rPAD/4791 PAD:6618 PAD:6619 1.5
rPAD/4792 PAD:6615 PAD:6618 0.0751765
rPAD/4793 PAD:6615 PAD:12323 1.5
rPAD/4794 PAD:6612 PAD:6615 0.0375882
rPAD/4795 PAD:6612 PAD:12320 1.5
rPAD/4796 PAD:6610 PAD:12320 0.0751765
rPAD/4797 PAD:6610 PAD:12318 1.5
rPAD/4798 PAD:6609 PAD:6612 0.0751765
rPAD/4799 PAD:6609 PAD:6610 1.5
rPAD/4800 PAD:6607 PAD:6610 0.0375882
rPAD/4801 PAD:6607 PAD:12315 1.5
rPAD/4802 PAD:6606 PAD:6609 0.0375882
rPAD/4803 PAD:6606 PAD:6607 1.5
rPAD/4804 PAD:6604 PAD:6607 0.0751765
rPAD/4805 PAD:6604 PAD:12312 1.5
rPAD/4806 PAD:6603 PAD:6606 0.0751765
rPAD/4807 PAD:6603 PAD:6604 1.5
rPAD/4808 PAD:6601 PAD:6604 0.0375882
rPAD/4809 PAD:6601 PAD:12309 1.5
rPAD/4810 PAD:6600 PAD:6603 0.0375882
rPAD/4811 PAD:6600 PAD:6601 1.5
rPAD/4812 PAD:6598 PAD:6601 0.0751765
rPAD/4813 PAD:6598 PAD:12306 1.5
rPAD/4814 PAD:6597 PAD:6600 0.0751765
rPAD/4815 PAD:6597 PAD:6598 1.5
rPAD/4816 PAD:6595 PAD:12299 0.0751765
rPAD/4817 PAD:6595 PAD:6598 0.0375882
rPAD/4818 PAD:6595 PAD:12303 1.5
rPAD/4819 PAD:6594 PAD:6597 0.0375882
rPAD/4820 PAD:6594 PAD:6595 1.5
rPAD/4821 PAD:6591 PAD:6594 0.0751765
rPAD/4822 PAD:6591 PAD:12299 1.5
rPAD/4823 PAD:6589 PAD:12299 0.0375882
rPAD/4824 PAD:6589 PAD:12297 1.5
rPAD/4825 PAD:6588 PAD:6591 0.0375882
rPAD/4826 PAD:6588 PAD:6589 1.5
rPAD/4827 PAD:6586 PAD:6589 0.0751765
rPAD/4828 PAD:6586 PAD:12294 1.5
rPAD/4829 PAD:6585 PAD:6588 0.0751765
rPAD/4830 PAD:6585 PAD:6586 1.5
rPAD/4831 PAD:6583 PAD:12287 0.0751765
rPAD/4832 PAD:6583 PAD:6586 0.0375882
rPAD/4833 PAD:6583 PAD:12291 1.5
rPAD/4834 PAD:6582 PAD:6585 0.0375882
rPAD/4835 PAD:6582 PAD:6583 1.5
rPAD/4836 PAD:6579 PAD:6582 0.0751765
rPAD/4837 PAD:6579 PAD:12287 1.5
rPAD/4838 PAD:6576 PAD:6579 0.0375882
rPAD/4839 PAD:6576 PAD:12284 1.5
rPAD/4840 PAD:6573 PAD:6576 0.0751765
rPAD/4841 PAD:6573 PAD:12281 1.5
rPAD/4842 PAD:6570 PAD:6573 0.0375882
rPAD/4843 PAD:6570 PAD:12278 1.5
rPAD/4844 PAD:6567 PAD:6570 0.0751765
rPAD/4845 PAD:6567 PAD:12275 1.5
rPAD/4846 PAD:6565 PAD:12275 0.0375882
rPAD/4847 PAD:6565 PAD:12273 1.5
rPAD/4848 PAD:6564 PAD:6567 0.0375882
rPAD/4849 PAD:6564 PAD:6565 1.5
rPAD/4850 PAD:6562 PAD:12266 0.0375882
rPAD/4851 PAD:6562 PAD:6565 0.0751765
rPAD/4852 PAD:6562 PAD:12270 1.5
rPAD/4853 PAD:6561 PAD:6564 0.0751765
rPAD/4854 PAD:6561 PAD:6562 1.5
rPAD/4855 PAD:6558 PAD:6561 0.0375882
rPAD/4856 PAD:6558 PAD:12266 1.5
rPAD/4857 PAD:6556 PAD:12266 0.0751765
rPAD/4858 PAD:6556 PAD:12264 1.5
rPAD/4859 PAD:6555 PAD:6558 0.0751765
rPAD/4860 PAD:6555 PAD:6556 1.5
rPAD/4861 PAD:6553 PAD:6556 0.0375882
rPAD/4862 PAD:6553 PAD:12261 1.5
rPAD/4863 PAD:6552 PAD:6555 0.0375882
rPAD/4864 PAD:6552 PAD:6553 1.5
rPAD/4865 PAD:6550 PAD:6553 0.0751765
rPAD/4866 PAD:6550 PAD:12258 1.5
rPAD/4867 PAD:6549 PAD:6552 0.0751765
rPAD/4868 PAD:6549 PAD:6550 1.5
rPAD/4869 PAD:6547 PAD:6550 0.0375882
rPAD/4870 PAD:6547 PAD:12255 1.5
rPAD/4871 PAD:6546 PAD:6549 0.0375882
rPAD/4872 PAD:6546 PAD:6547 1.5
rPAD/4873 PAD:6544 PAD:6547 0.0751765
rPAD/4874 PAD:6544 PAD:12252 1.5
rPAD/4875 PAD:6543 PAD:6546 0.0751765
rPAD/4876 PAD:6543 PAD:6544 1.5
rPAD/4877 PAD:6541 PAD:12245 0.0751765
rPAD/4878 PAD:6541 PAD:6544 0.0375882
rPAD/4879 PAD:6541 PAD:12249 1.5
rPAD/4880 PAD:6540 PAD:6543 0.0375882
rPAD/4881 PAD:6540 PAD:6541 1.5
rPAD/4882 PAD:6537 PAD:6540 0.0751765
rPAD/4883 PAD:6537 PAD:12245 1.5
rPAD/4884 PAD:6535 PAD:12245 0.0375882
rPAD/4885 PAD:6535 PAD:12243 1.5
rPAD/4886 PAD:6534 PAD:6537 0.0375882
rPAD/4887 PAD:6534 PAD:6535 1.5
rPAD/4888 PAD:6532 PAD:6535 0.0751765
rPAD/4889 PAD:6532 PAD:12240 1.5
rPAD/4890 PAD:6531 PAD:6534 0.0751765
rPAD/4891 PAD:6531 PAD:6532 1.5
rPAD/4892 PAD:6529 PAD:6532 0.0375882
rPAD/4893 PAD:6529 PAD:12237 1.5
rPAD/4894 PAD:6528 PAD:6531 0.0375882
rPAD/4895 PAD:6528 PAD:6529 1.5
rPAD/4896 PAD:6526 PAD:6529 0.0751765
rPAD/4897 PAD:6526 PAD:12234 1.5
rPAD/4898 PAD:6525 PAD:6528 0.0751765
rPAD/4899 PAD:6525 PAD:6526 1.5
rPAD/4900 PAD:6523 PAD:6526 0.0375882
rPAD/4901 PAD:6523 PAD:12231 1.5
rPAD/4902 PAD:6522 PAD:6525 0.0375882
rPAD/4903 PAD:6522 PAD:6523 1.5
rPAD/4904 PAD:6520 PAD:6523 0.0751765
rPAD/4905 PAD:6520 PAD:12228 1.5
rPAD/4906 PAD:6519 PAD:6522 0.0751765
rPAD/4907 PAD:6519 PAD:6520 1.5
rPAD/4908 PAD:6517 PAD:6520 0.0375882
rPAD/4909 PAD:6517 PAD:12225 1.5
rPAD/4910 PAD:6516 PAD:6519 0.0375882
rPAD/4911 PAD:6516 PAD:6517 1.5
rPAD/4912 PAD:6514 PAD:14916 0.0283817
rPAD/4913 PAD:6514 PAD:6517 0.0751765
rPAD/4914 PAD:6514 PAD:12222 1.5
rPAD/4915 PAD:6513 PAD:9203 0.0378785
rPAD/4916 PAD:6513 PAD:6516 0.0751765
rPAD/4917 PAD:6513 PAD:6514 1.5
rPAD/4918 PAD:6509 PAD:12049 0.0100588
rPAD/4919 PAD:6509 PAD:12217 1.5
rPAD/4920 PAD:6508 PAD:9379 0.0670908
rPAD/4921 PAD:6508 PAD:6509 1.5
rPAD/4922 PAD:6506 PAD:6509 0.0751765
rPAD/4923 PAD:6506 PAD:12214 1.5
rPAD/4924 PAD:6505 PAD:6508 0.0751765
rPAD/4925 PAD:6505 PAD:6506 1.5
rPAD/4926 PAD:6503 PAD:12207 0.0751765
rPAD/4927 PAD:6503 PAD:6506 0.0375882
rPAD/4928 PAD:6503 PAD:12211 1.5
rPAD/4929 PAD:6502 PAD:6505 0.0375882
rPAD/4930 PAD:6502 PAD:6503 1.5
rPAD/4931 PAD:6499 PAD:6502 0.0751765
rPAD/4932 PAD:6499 PAD:12207 1.5
rPAD/4933 PAD:6497 PAD:12207 0.0375882
rPAD/4934 PAD:6497 PAD:12205 1.5
rPAD/4935 PAD:6496 PAD:6499 0.0375882
rPAD/4936 PAD:6496 PAD:6497 1.5
rPAD/4937 PAD:6494 PAD:6497 0.0751765
rPAD/4938 PAD:6494 PAD:12202 1.5
rPAD/4939 PAD:6493 PAD:6496 0.0751765
rPAD/4940 PAD:6493 PAD:6494 1.5
rPAD/4941 PAD:6491 PAD:6494 0.0375882
rPAD/4942 PAD:6491 PAD:12199 1.5
rPAD/4943 PAD:6490 PAD:6493 0.0375882
rPAD/4944 PAD:6490 PAD:6491 1.5
rPAD/4945 PAD:6488 PAD:6491 0.0751765
rPAD/4946 PAD:6488 PAD:12196 1.5
rPAD/4947 PAD:6487 PAD:6490 0.0751765
rPAD/4948 PAD:6487 PAD:6488 1.5
rPAD/4949 PAD:6485 PAD:6488 0.0375882
rPAD/4950 PAD:6485 PAD:12193 1.5
rPAD/4951 PAD:6484 PAD:6487 0.0375882
rPAD/4952 PAD:6484 PAD:6485 1.5
rPAD/4953 PAD:6482 PAD:6485 0.0751765
rPAD/4954 PAD:6482 PAD:12190 1.5
rPAD/4955 PAD:6481 PAD:6484 0.0751765
rPAD/4956 PAD:6481 PAD:6482 1.5
rPAD/4957 PAD:6479 PAD:6482 0.0375882
rPAD/4958 PAD:6479 PAD:12187 1.5
rPAD/4959 PAD:6478 PAD:6481 0.0375882
rPAD/4960 PAD:6478 PAD:6479 1.5
rPAD/4961 PAD:6476 PAD:6479 0.0751765
rPAD/4962 PAD:6476 PAD:12184 1.5
rPAD/4963 PAD:6475 PAD:6478 0.0751765
rPAD/4964 PAD:6475 PAD:6476 1.5
rPAD/4965 PAD:6473 PAD:6476 0.0375882
rPAD/4966 PAD:6473 PAD:12181 1.5
rPAD/4967 PAD:6472 PAD:6475 0.0375882
rPAD/4968 PAD:6472 PAD:6473 1.5
rPAD/4969 PAD:6470 PAD:6473 0.0751765
rPAD/4970 PAD:6470 PAD:12178 1.5
rPAD/4971 PAD:6469 PAD:6472 0.0751765
rPAD/4972 PAD:6469 PAD:6470 1.5
rPAD/4973 PAD:6467 PAD:12171 0.0751765
rPAD/4974 PAD:6467 PAD:6470 0.0375882
rPAD/4975 PAD:6467 PAD:12175 1.5
rPAD/4976 PAD:6466 PAD:6469 0.0375882
rPAD/4977 PAD:6466 PAD:6467 1.5
rPAD/4978 PAD:6463 PAD:6466 0.0751765
rPAD/4979 PAD:6463 PAD:12171 1.5
rPAD/4980 PAD:6461 PAD:12165 0.0751765
rPAD/4981 PAD:6461 PAD:12171 0.0375882
rPAD/4982 PAD:6461 PAD:12169 1.5
rPAD/4983 PAD:6460 PAD:6463 0.0375882
rPAD/4984 PAD:6460 PAD:6461 1.5
rPAD/4985 PAD:6457 PAD:6460 0.0751765
rPAD/4986 PAD:6457 PAD:12165 1.5
rPAD/4987 PAD:6454 PAD:6457 0.0375882
rPAD/4988 PAD:6454 PAD:12162 1.5
rPAD/4989 PAD:6451 PAD:6454 0.0751765
rPAD/4990 PAD:6451 PAD:12159 1.5
rPAD/4991 PAD:6449 PAD:12153 0.0751765
rPAD/4992 PAD:6449 PAD:12159 0.0375882
rPAD/4993 PAD:6449 PAD:12157 1.5
rPAD/4994 PAD:6448 PAD:6451 0.0375882
rPAD/4995 PAD:6448 PAD:6449 1.5
rPAD/4996 PAD:6445 PAD:6448 0.0751765
rPAD/4997 PAD:6445 PAD:12153 1.5
rPAD/4998 PAD:6442 PAD:6445 0.0375882
rPAD/4999 PAD:6442 PAD:12150 1.5
rPAD/5000 PAD:6440 PAD:12150 0.0751765
rPAD/5001 PAD:6440 PAD:12148 1.5
rPAD/5002 PAD:6439 PAD:6442 0.0751765
rPAD/5003 PAD:6439 PAD:6440 1.5
rPAD/5004 PAD:6437 PAD:6440 0.0375882
rPAD/5005 PAD:6437 PAD:12145 1.5
rPAD/5006 PAD:6436 PAD:6439 0.0375882
rPAD/5007 PAD:6436 PAD:6437 1.5
rPAD/5008 PAD:6434 PAD:6437 0.0751765
rPAD/5009 PAD:6434 PAD:12142 1.5
rPAD/5010 PAD:6433 PAD:6436 0.0751765
rPAD/5011 PAD:6433 PAD:6434 1.5
rPAD/5012 PAD:6431 PAD:6434 0.0375882
rPAD/5013 PAD:6431 PAD:12139 1.5
rPAD/5014 PAD:6430 PAD:6433 0.0375882
rPAD/5015 PAD:6430 PAD:6431 1.5
rPAD/5016 PAD:6428 PAD:6431 0.0751765
rPAD/5017 PAD:6428 PAD:12136 1.5
rPAD/5018 PAD:6427 PAD:6430 0.0751765
rPAD/5019 PAD:6427 PAD:6428 1.5
rPAD/5020 PAD:6425 PAD:12129 0.0751765
rPAD/5021 PAD:6425 PAD:6428 0.0375882
rPAD/5022 PAD:6425 PAD:12133 1.5
rPAD/5023 PAD:6424 PAD:6427 0.0375882
rPAD/5024 PAD:6424 PAD:6425 1.5
rPAD/5025 PAD:6421 PAD:6424 0.0751765
rPAD/5026 PAD:6421 PAD:12129 1.5
rPAD/5027 PAD:6419 PAD:12129 0.0375882
rPAD/5028 PAD:6419 PAD:12127 1.5
rPAD/5029 PAD:6418 PAD:6421 0.0375882
rPAD/5030 PAD:6418 PAD:6419 1.5
rPAD/5031 PAD:6416 PAD:6419 0.0751765
rPAD/5032 PAD:6416 PAD:12124 1.5
rPAD/5033 PAD:6415 PAD:6418 0.0751765
rPAD/5034 PAD:6415 PAD:6416 1.5
rPAD/5035 PAD:6413 PAD:12117 0.0751765
rPAD/5036 PAD:6413 PAD:6416 0.0375882
rPAD/5037 PAD:6413 PAD:12121 1.5
rPAD/5038 PAD:6412 PAD:6415 0.0375882
rPAD/5039 PAD:6412 PAD:6413 1.5
rPAD/5040 PAD:6409 PAD:6412 0.0751765
rPAD/5041 PAD:6409 PAD:12117 1.5
rPAD/5042 PAD:6406 PAD:6409 0.0375882
rPAD/5043 PAD:6406 PAD:12114 1.5
rPAD/5044 PAD:6403 PAD:6406 0.0751765
rPAD/5045 PAD:6403 PAD:12111 1.5
rPAD/5046 PAD:6400 PAD:6403 0.0375882
rPAD/5047 PAD:6400 PAD:12108 1.5
rPAD/5048 PAD:6397 PAD:6400 0.0751765
rPAD/5049 PAD:6397 PAD:12105 1.5
rPAD/5050 PAD:6395 PAD:12105 0.0375882
rPAD/5051 PAD:6395 PAD:12103 1.5
rPAD/5052 PAD:6394 PAD:6397 0.0375882
rPAD/5053 PAD:6394 PAD:6395 1.5
rPAD/5054 PAD:6392 PAD:12096 0.0375882
rPAD/5055 PAD:6392 PAD:6395 0.0751765
rPAD/5056 PAD:6392 PAD:12100 1.5
rPAD/5057 PAD:6391 PAD:6394 0.0751765
rPAD/5058 PAD:6391 PAD:6392 1.5
rPAD/5059 PAD:6388 PAD:6391 0.0375882
rPAD/5060 PAD:6388 PAD:12096 1.5
rPAD/5061 PAD:6386 PAD:12096 0.0751765
rPAD/5062 PAD:6386 PAD:12094 1.5
rPAD/5063 PAD:6385 PAD:6388 0.0751765
rPAD/5064 PAD:6385 PAD:6386 1.5
rPAD/5065 PAD:6383 PAD:6386 0.0375882
rPAD/5066 PAD:6383 PAD:12091 1.5
rPAD/5067 PAD:6382 PAD:6385 0.0375882
rPAD/5068 PAD:6382 PAD:6383 1.5
rPAD/5069 PAD:6380 PAD:6383 0.0751765
rPAD/5070 PAD:6380 PAD:12088 1.5
rPAD/5071 PAD:6379 PAD:6382 0.0751765
rPAD/5072 PAD:6379 PAD:6380 1.5
rPAD/5073 PAD:6377 PAD:6380 0.0375882
rPAD/5074 PAD:6377 PAD:12085 1.5
rPAD/5075 PAD:6376 PAD:6379 0.0375882
rPAD/5076 PAD:6376 PAD:6377 1.5
rPAD/5077 PAD:6374 PAD:6377 0.0751765
rPAD/5078 PAD:6374 PAD:12082 1.5
rPAD/5079 PAD:6373 PAD:6376 0.0751765
rPAD/5080 PAD:6373 PAD:6374 1.5
rPAD/5081 PAD:6371 PAD:12075 0.0751765
rPAD/5082 PAD:6371 PAD:6374 0.0375882
rPAD/5083 PAD:6371 PAD:12079 1.5
rPAD/5084 PAD:6370 PAD:6373 0.0375882
rPAD/5085 PAD:6370 PAD:6371 1.5
rPAD/5086 PAD:6367 PAD:6370 0.0751765
rPAD/5087 PAD:6367 PAD:12075 1.5
rPAD/5088 PAD:6365 PAD:12075 0.0375882
rPAD/5089 PAD:6365 PAD:12073 1.5
rPAD/5090 PAD:6364 PAD:6367 0.0375882
rPAD/5091 PAD:6364 PAD:6365 1.5
rPAD/5092 PAD:6362 PAD:6365 0.0751765
rPAD/5093 PAD:6362 PAD:12070 1.5
rPAD/5094 PAD:6361 PAD:6364 0.0751765
rPAD/5095 PAD:6361 PAD:6362 1.5
rPAD/5096 PAD:6359 PAD:6362 0.0375882
rPAD/5097 PAD:6359 PAD:12067 1.5
rPAD/5098 PAD:6358 PAD:6361 0.0375882
rPAD/5099 PAD:6358 PAD:6359 1.5
rPAD/5100 PAD:6356 PAD:6359 0.0751765
rPAD/5101 PAD:6356 PAD:12064 1.5
rPAD/5102 PAD:6355 PAD:6358 0.0751765
rPAD/5103 PAD:6355 PAD:6356 1.5
rPAD/5104 PAD:6353 PAD:6356 0.0375882
rPAD/5105 PAD:6353 PAD:12061 1.5
rPAD/5106 PAD:6352 PAD:6355 0.0375882
rPAD/5107 PAD:6352 PAD:6353 1.5
rPAD/5108 PAD:6350 PAD:6353 0.0751765
rPAD/5109 PAD:6350 PAD:12058 1.5
rPAD/5110 PAD:6349 PAD:6352 0.0751765
rPAD/5111 PAD:6349 PAD:6350 1.5
rPAD/5112 PAD:6347 PAD:6350 0.0375882
rPAD/5113 PAD:6347 PAD:12055 1.5
rPAD/5114 PAD:6346 PAD:6349 0.0375882
rPAD/5115 PAD:6346 PAD:6347 1.5
rPAD/5116 PAD:6344 PAD:14911 0.0283817
rPAD/5117 PAD:6344 PAD:6347 0.0751765
rPAD/5118 PAD:6344 PAD:12052 1.5
rPAD/5119 PAD:6343 PAD:9196 0.0378785
rPAD/5120 PAD:6343 PAD:6346 0.0751765
rPAD/5121 PAD:6343 PAD:6344 1.5
rPAD/5122 PAD:6339 PAD:11879 0.0100588
rPAD/5123 PAD:6339 PAD:12047 1.5
rPAD/5124 PAD:6338 PAD:9375 0.0670908
rPAD/5125 PAD:6338 PAD:6339 1.5
rPAD/5126 PAD:6336 PAD:6339 0.0751765
rPAD/5127 PAD:6336 PAD:12044 1.5
rPAD/5128 PAD:6335 PAD:6338 0.0751765
rPAD/5129 PAD:6335 PAD:6336 1.5
rPAD/5130 PAD:6333 PAD:12037 0.0751765
rPAD/5131 PAD:6333 PAD:6336 0.0375882
rPAD/5132 PAD:6333 PAD:12041 1.5
rPAD/5133 PAD:6332 PAD:6335 0.0375882
rPAD/5134 PAD:6332 PAD:6333 1.5
rPAD/5135 PAD:6329 PAD:6332 0.0751765
rPAD/5136 PAD:6329 PAD:12037 1.5
rPAD/5137 PAD:6327 PAD:12037 0.0375882
rPAD/5138 PAD:6327 PAD:12035 1.5
rPAD/5139 PAD:6326 PAD:6329 0.0375882
rPAD/5140 PAD:6326 PAD:6327 1.5
rPAD/5141 PAD:6324 PAD:6327 0.0751765
rPAD/5142 PAD:6324 PAD:12032 1.5
rPAD/5143 PAD:6323 PAD:6326 0.0751765
rPAD/5144 PAD:6323 PAD:6324 1.5
rPAD/5145 PAD:6321 PAD:6324 0.0375882
rPAD/5146 PAD:6321 PAD:12029 1.5
rPAD/5147 PAD:6320 PAD:6323 0.0375882
rPAD/5148 PAD:6320 PAD:6321 1.5
rPAD/5149 PAD:6318 PAD:6321 0.0751765
rPAD/5150 PAD:6318 PAD:12026 1.5
rPAD/5151 PAD:6317 PAD:6320 0.0751765
rPAD/5152 PAD:6317 PAD:6318 1.5
rPAD/5153 PAD:6315 PAD:6318 0.0375882
rPAD/5154 PAD:6315 PAD:12023 1.5
rPAD/5155 PAD:6314 PAD:6317 0.0375882
rPAD/5156 PAD:6314 PAD:6315 1.5
rPAD/5157 PAD:6312 PAD:6315 0.0751765
rPAD/5158 PAD:6312 PAD:12020 1.5
rPAD/5159 PAD:6311 PAD:6314 0.0751765
rPAD/5160 PAD:6311 PAD:6312 1.5
rPAD/5161 PAD:6309 PAD:6312 0.0375882
rPAD/5162 PAD:6309 PAD:12017 1.5
rPAD/5163 PAD:6308 PAD:6311 0.0375882
rPAD/5164 PAD:6308 PAD:6309 1.5
rPAD/5165 PAD:6306 PAD:6309 0.0751765
rPAD/5166 PAD:6306 PAD:12014 1.5
rPAD/5167 PAD:6305 PAD:6308 0.0751765
rPAD/5168 PAD:6305 PAD:6306 1.5
rPAD/5169 PAD:6303 PAD:6306 0.0375882
rPAD/5170 PAD:6303 PAD:12011 1.5
rPAD/5171 PAD:6302 PAD:6305 0.0375882
rPAD/5172 PAD:6302 PAD:6303 1.5
rPAD/5173 PAD:6300 PAD:6303 0.0751765
rPAD/5174 PAD:6300 PAD:12008 1.5
rPAD/5175 PAD:6299 PAD:6302 0.0751765
rPAD/5176 PAD:6299 PAD:6300 1.5
rPAD/5177 PAD:6297 PAD:12001 0.0751765
rPAD/5178 PAD:6297 PAD:6300 0.0375882
rPAD/5179 PAD:6297 PAD:12005 1.5
rPAD/5180 PAD:6296 PAD:6299 0.0375882
rPAD/5181 PAD:6296 PAD:6297 1.5
rPAD/5182 PAD:6293 PAD:6296 0.0751765
rPAD/5183 PAD:6293 PAD:12001 1.5
rPAD/5184 PAD:6291 PAD:11995 0.0751765
rPAD/5185 PAD:6291 PAD:12001 0.0375882
rPAD/5186 PAD:6291 PAD:11999 1.5
rPAD/5187 PAD:6290 PAD:6293 0.0375882
rPAD/5188 PAD:6290 PAD:6291 1.5
rPAD/5189 PAD:6287 PAD:6290 0.0751765
rPAD/5190 PAD:6287 PAD:11995 1.5
rPAD/5191 PAD:6284 PAD:6287 0.0375882
rPAD/5192 PAD:6284 PAD:11992 1.5
rPAD/5193 PAD:6281 PAD:6284 0.0751765
rPAD/5194 PAD:6281 PAD:11989 1.5
rPAD/5195 PAD:6279 PAD:11983 0.0751765
rPAD/5196 PAD:6279 PAD:11989 0.0375882
rPAD/5197 PAD:6279 PAD:11987 1.5
rPAD/5198 PAD:6278 PAD:6281 0.0375882
rPAD/5199 PAD:6278 PAD:6279 1.5
rPAD/5200 PAD:6275 PAD:6278 0.0751765
rPAD/5201 PAD:6275 PAD:11983 1.5
rPAD/5202 PAD:6272 PAD:6275 0.0375882
rPAD/5203 PAD:6272 PAD:11980 1.5
rPAD/5204 PAD:6270 PAD:11980 0.0751765
rPAD/5205 PAD:6270 PAD:11978 1.5
rPAD/5206 PAD:6269 PAD:6272 0.0751765
rPAD/5207 PAD:6269 PAD:6270 1.5
rPAD/5208 PAD:6267 PAD:6270 0.0375882
rPAD/5209 PAD:6267 PAD:11975 1.5
rPAD/5210 PAD:6266 PAD:6269 0.0375882
rPAD/5211 PAD:6266 PAD:6267 1.5
rPAD/5212 PAD:6264 PAD:6267 0.0751765
rPAD/5213 PAD:6264 PAD:11972 1.5
rPAD/5214 PAD:6263 PAD:6266 0.0751765
rPAD/5215 PAD:6263 PAD:6264 1.5
rPAD/5216 PAD:6261 PAD:6264 0.0375882
rPAD/5217 PAD:6261 PAD:11969 1.5
rPAD/5218 PAD:6260 PAD:6263 0.0375882
rPAD/5219 PAD:6260 PAD:6261 1.5
rPAD/5220 PAD:6258 PAD:6261 0.0751765
rPAD/5221 PAD:6258 PAD:11966 1.5
rPAD/5222 PAD:6257 PAD:6260 0.0751765
rPAD/5223 PAD:6257 PAD:6258 1.5
rPAD/5224 PAD:6255 PAD:11959 0.0751765
rPAD/5225 PAD:6255 PAD:6258 0.0375882
rPAD/5226 PAD:6255 PAD:11963 1.5
rPAD/5227 PAD:6254 PAD:6257 0.0375882
rPAD/5228 PAD:6254 PAD:6255 1.5
rPAD/5229 PAD:6251 PAD:6254 0.0751765
rPAD/5230 PAD:6251 PAD:11959 1.5
rPAD/5231 PAD:6249 PAD:11959 0.0375882
rPAD/5232 PAD:6249 PAD:11957 1.5
rPAD/5233 PAD:6248 PAD:6251 0.0375882
rPAD/5234 PAD:6248 PAD:6249 1.5
rPAD/5235 PAD:6246 PAD:6249 0.0751765
rPAD/5236 PAD:6246 PAD:11954 1.5
rPAD/5237 PAD:6245 PAD:6248 0.0751765
rPAD/5238 PAD:6245 PAD:6246 1.5
rPAD/5239 PAD:6243 PAD:11947 0.0751765
rPAD/5240 PAD:6243 PAD:6246 0.0375882
rPAD/5241 PAD:6243 PAD:11951 1.5
rPAD/5242 PAD:6242 PAD:6245 0.0375882
rPAD/5243 PAD:6242 PAD:6243 1.5
rPAD/5244 PAD:6239 PAD:6242 0.0751765
rPAD/5245 PAD:6239 PAD:11947 1.5
rPAD/5246 PAD:6236 PAD:6239 0.0375882
rPAD/5247 PAD:6236 PAD:11944 1.5
rPAD/5248 PAD:6233 PAD:6236 0.0751765
rPAD/5249 PAD:6233 PAD:11941 1.5
rPAD/5250 PAD:6230 PAD:6233 0.0375882
rPAD/5251 PAD:6230 PAD:11938 1.5
rPAD/5252 PAD:6227 PAD:6230 0.0751765
rPAD/5253 PAD:6227 PAD:11935 1.5
rPAD/5254 PAD:6225 PAD:11935 0.0375882
rPAD/5255 PAD:6225 PAD:11933 1.5
rPAD/5256 PAD:6224 PAD:6227 0.0375882
rPAD/5257 PAD:6224 PAD:6225 1.5
rPAD/5258 PAD:6222 PAD:11926 0.0375882
rPAD/5259 PAD:6222 PAD:6225 0.0751765
rPAD/5260 PAD:6222 PAD:11930 1.5
rPAD/5261 PAD:6221 PAD:6224 0.0751765
rPAD/5262 PAD:6221 PAD:6222 1.5
rPAD/5263 PAD:6218 PAD:6221 0.0375882
rPAD/5264 PAD:6218 PAD:11926 1.5
rPAD/5265 PAD:6216 PAD:11926 0.0751765
rPAD/5266 PAD:6216 PAD:11924 1.5
rPAD/5267 PAD:6215 PAD:6218 0.0751765
rPAD/5268 PAD:6215 PAD:6216 1.5
rPAD/5269 PAD:6213 PAD:6216 0.0375882
rPAD/5270 PAD:6213 PAD:11921 1.5
rPAD/5271 PAD:6212 PAD:6215 0.0375882
rPAD/5272 PAD:6212 PAD:6213 1.5
rPAD/5273 PAD:6210 PAD:6213 0.0751765
rPAD/5274 PAD:6210 PAD:11918 1.5
rPAD/5275 PAD:6209 PAD:6212 0.0751765
rPAD/5276 PAD:6209 PAD:6210 1.5
rPAD/5277 PAD:6207 PAD:6210 0.0375882
rPAD/5278 PAD:6207 PAD:11915 1.5
rPAD/5279 PAD:6206 PAD:6209 0.0375882
rPAD/5280 PAD:6206 PAD:6207 1.5
rPAD/5281 PAD:6204 PAD:6207 0.0751765
rPAD/5282 PAD:6204 PAD:11912 1.5
rPAD/5283 PAD:6203 PAD:6206 0.0751765
rPAD/5284 PAD:6203 PAD:6204 1.5
rPAD/5285 PAD:6201 PAD:11905 0.0751765
rPAD/5286 PAD:6201 PAD:6204 0.0375882
rPAD/5287 PAD:6201 PAD:11909 1.5
rPAD/5288 PAD:6200 PAD:6203 0.0375882
rPAD/5289 PAD:6200 PAD:6201 1.5
rPAD/5290 PAD:6197 PAD:6200 0.0751765
rPAD/5291 PAD:6197 PAD:11905 1.5
rPAD/5292 PAD:6195 PAD:11905 0.0375882
rPAD/5293 PAD:6195 PAD:11903 1.5
rPAD/5294 PAD:6194 PAD:6197 0.0375882
rPAD/5295 PAD:6194 PAD:6195 1.5
rPAD/5296 PAD:6192 PAD:6195 0.0751765
rPAD/5297 PAD:6192 PAD:11900 1.5
rPAD/5298 PAD:6191 PAD:6194 0.0751765
rPAD/5299 PAD:6191 PAD:6192 1.5
rPAD/5300 PAD:6189 PAD:6192 0.0375882
rPAD/5301 PAD:6189 PAD:11897 1.5
rPAD/5302 PAD:6188 PAD:6191 0.0375882
rPAD/5303 PAD:6188 PAD:6189 1.5
rPAD/5304 PAD:6186 PAD:6189 0.0751765
rPAD/5305 PAD:6186 PAD:11894 1.5
rPAD/5306 PAD:6185 PAD:6188 0.0751765
rPAD/5307 PAD:6185 PAD:6186 1.5
rPAD/5308 PAD:6183 PAD:6186 0.0375882
rPAD/5309 PAD:6183 PAD:11891 1.5
rPAD/5310 PAD:6182 PAD:6185 0.0375882
rPAD/5311 PAD:6182 PAD:6183 1.5
rPAD/5312 PAD:6180 PAD:6183 0.0751765
rPAD/5313 PAD:6180 PAD:11888 1.5
rPAD/5314 PAD:6179 PAD:6182 0.0751765
rPAD/5315 PAD:6179 PAD:6180 1.5
rPAD/5316 PAD:6177 PAD:6180 0.0375882
rPAD/5317 PAD:6177 PAD:11885 1.5
rPAD/5318 PAD:6176 PAD:6179 0.0375882
rPAD/5319 PAD:6176 PAD:6177 1.5
rPAD/5320 PAD:6174 PAD:14906 0.0283817
rPAD/5321 PAD:6174 PAD:6177 0.0751765
rPAD/5322 PAD:6174 PAD:11882 1.5
rPAD/5323 PAD:6173 PAD:9189 0.0378785
rPAD/5324 PAD:6173 PAD:6176 0.0751765
rPAD/5325 PAD:6173 PAD:6174 1.5
rPAD/5326 PAD:6169 PAD:11709 0.0100588
rPAD/5327 PAD:6169 PAD:11877 1.5
rPAD/5328 PAD:6168 PAD:9371 0.0670908
rPAD/5329 PAD:6168 PAD:6169 1.5
rPAD/5330 PAD:6166 PAD:6169 0.0751765
rPAD/5331 PAD:6166 PAD:11874 1.5
rPAD/5332 PAD:6165 PAD:6168 0.0751765
rPAD/5333 PAD:6165 PAD:6166 1.5
rPAD/5334 PAD:6163 PAD:11867 0.0751765
rPAD/5335 PAD:6163 PAD:6166 0.0375882
rPAD/5336 PAD:6163 PAD:11871 1.5
rPAD/5337 PAD:6162 PAD:6165 0.0375882
rPAD/5338 PAD:6162 PAD:6163 1.5
rPAD/5339 PAD:6159 PAD:6162 0.0751765
rPAD/5340 PAD:6159 PAD:11867 1.5
rPAD/5341 PAD:6157 PAD:11867 0.0375882
rPAD/5342 PAD:6157 PAD:11865 1.5
rPAD/5343 PAD:6156 PAD:6159 0.0375882
rPAD/5344 PAD:6156 PAD:6157 1.5
rPAD/5345 PAD:6154 PAD:6157 0.0751765
rPAD/5346 PAD:6154 PAD:11862 1.5
rPAD/5347 PAD:6153 PAD:6156 0.0751765
rPAD/5348 PAD:6153 PAD:6154 1.5
rPAD/5349 PAD:6151 PAD:6154 0.0375882
rPAD/5350 PAD:6151 PAD:11859 1.5
rPAD/5351 PAD:6150 PAD:6153 0.0375882
rPAD/5352 PAD:6150 PAD:6151 1.5
rPAD/5353 PAD:6148 PAD:6151 0.0751765
rPAD/5354 PAD:6148 PAD:11856 1.5
rPAD/5355 PAD:6147 PAD:6150 0.0751765
rPAD/5356 PAD:6147 PAD:6148 1.5
rPAD/5357 PAD:6145 PAD:6148 0.0375882
rPAD/5358 PAD:6145 PAD:11853 1.5
rPAD/5359 PAD:6144 PAD:6147 0.0375882
rPAD/5360 PAD:6144 PAD:6145 1.5
rPAD/5361 PAD:6142 PAD:6145 0.0751765
rPAD/5362 PAD:6142 PAD:11850 1.5
rPAD/5363 PAD:6141 PAD:6144 0.0751765
rPAD/5364 PAD:6141 PAD:6142 1.5
rPAD/5365 PAD:6139 PAD:6142 0.0375882
rPAD/5366 PAD:6139 PAD:11847 1.5
rPAD/5367 PAD:6138 PAD:6141 0.0375882
rPAD/5368 PAD:6138 PAD:6139 1.5
rPAD/5369 PAD:6136 PAD:6139 0.0751765
rPAD/5370 PAD:6136 PAD:11844 1.5
rPAD/5371 PAD:6135 PAD:6138 0.0751765
rPAD/5372 PAD:6135 PAD:6136 1.5
rPAD/5373 PAD:6133 PAD:6136 0.0375882
rPAD/5374 PAD:6133 PAD:11841 1.5
rPAD/5375 PAD:6132 PAD:6135 0.0375882
rPAD/5376 PAD:6132 PAD:6133 1.5
rPAD/5377 PAD:6130 PAD:6133 0.0751765
rPAD/5378 PAD:6130 PAD:11838 1.5
rPAD/5379 PAD:6129 PAD:6132 0.0751765
rPAD/5380 PAD:6129 PAD:6130 1.5
rPAD/5381 PAD:6127 PAD:11831 0.0751765
rPAD/5382 PAD:6127 PAD:6130 0.0375882
rPAD/5383 PAD:6127 PAD:11835 1.5
rPAD/5384 PAD:6126 PAD:6129 0.0375882
rPAD/5385 PAD:6126 PAD:6127 1.5
rPAD/5386 PAD:6123 PAD:6126 0.0751765
rPAD/5387 PAD:6123 PAD:11831 1.5
rPAD/5388 PAD:6121 PAD:11825 0.0751765
rPAD/5389 PAD:6121 PAD:11831 0.0375882
rPAD/5390 PAD:6121 PAD:11829 1.5
rPAD/5391 PAD:6120 PAD:6123 0.0375882
rPAD/5392 PAD:6120 PAD:6121 1.5
rPAD/5393 PAD:6117 PAD:6120 0.0751765
rPAD/5394 PAD:6117 PAD:11825 1.5
rPAD/5395 PAD:6114 PAD:6117 0.0375882
rPAD/5396 PAD:6114 PAD:11822 1.5
rPAD/5397 PAD:6111 PAD:6114 0.0751765
rPAD/5398 PAD:6111 PAD:11819 1.5
rPAD/5399 PAD:6109 PAD:11813 0.0751765
rPAD/5400 PAD:6109 PAD:11819 0.0375882
rPAD/5401 PAD:6109 PAD:11817 1.5
rPAD/5402 PAD:6108 PAD:6111 0.0375882
rPAD/5403 PAD:6108 PAD:6109 1.5
rPAD/5404 PAD:6105 PAD:6108 0.0751765
rPAD/5405 PAD:6105 PAD:11813 1.5
rPAD/5406 PAD:6102 PAD:6105 0.0375882
rPAD/5407 PAD:6102 PAD:11810 1.5
rPAD/5408 PAD:6100 PAD:11810 0.0751765
rPAD/5409 PAD:6100 PAD:11808 1.5
rPAD/5410 PAD:6099 PAD:6102 0.0751765
rPAD/5411 PAD:6099 PAD:6100 1.5
rPAD/5412 PAD:6097 PAD:6100 0.0375882
rPAD/5413 PAD:6097 PAD:11805 1.5
rPAD/5414 PAD:6096 PAD:6099 0.0375882
rPAD/5415 PAD:6096 PAD:6097 1.5
rPAD/5416 PAD:6094 PAD:6097 0.0751765
rPAD/5417 PAD:6094 PAD:11802 1.5
rPAD/5418 PAD:6093 PAD:6096 0.0751765
rPAD/5419 PAD:6093 PAD:6094 1.5
rPAD/5420 PAD:6091 PAD:6094 0.0375882
rPAD/5421 PAD:6091 PAD:11799 1.5
rPAD/5422 PAD:6090 PAD:6093 0.0375882
rPAD/5423 PAD:6090 PAD:6091 1.5
rPAD/5424 PAD:6088 PAD:6091 0.0751765
rPAD/5425 PAD:6088 PAD:11796 1.5
rPAD/5426 PAD:6087 PAD:6090 0.0751765
rPAD/5427 PAD:6087 PAD:6088 1.5
rPAD/5428 PAD:6085 PAD:11789 0.0751765
rPAD/5429 PAD:6085 PAD:6088 0.0375882
rPAD/5430 PAD:6085 PAD:11793 1.5
rPAD/5431 PAD:6084 PAD:6087 0.0375882
rPAD/5432 PAD:6084 PAD:6085 1.5
rPAD/5433 PAD:6081 PAD:6084 0.0751765
rPAD/5434 PAD:6081 PAD:11789 1.5
rPAD/5435 PAD:6079 PAD:11789 0.0375882
rPAD/5436 PAD:6079 PAD:11787 1.5
rPAD/5437 PAD:6078 PAD:6081 0.0375882
rPAD/5438 PAD:6078 PAD:6079 1.5
rPAD/5439 PAD:6076 PAD:6079 0.0751765
rPAD/5440 PAD:6076 PAD:11784 1.5
rPAD/5441 PAD:6075 PAD:6078 0.0751765
rPAD/5442 PAD:6075 PAD:6076 1.5
rPAD/5443 PAD:6073 PAD:11777 0.0751765
rPAD/5444 PAD:6073 PAD:6076 0.0375882
rPAD/5445 PAD:6073 PAD:11781 1.5
rPAD/5446 PAD:6072 PAD:6075 0.0375882
rPAD/5447 PAD:6072 PAD:6073 1.5
rPAD/5448 PAD:6069 PAD:6072 0.0751765
rPAD/5449 PAD:6069 PAD:11777 1.5
rPAD/5450 PAD:6066 PAD:6069 0.0375882
rPAD/5451 PAD:6066 PAD:11774 1.5
rPAD/5452 PAD:6063 PAD:6066 0.0751765
rPAD/5453 PAD:6063 PAD:11771 1.5
rPAD/5454 PAD:6060 PAD:6063 0.0375882
rPAD/5455 PAD:6060 PAD:11768 1.5
rPAD/5456 PAD:6057 PAD:6060 0.0751765
rPAD/5457 PAD:6057 PAD:11765 1.5
rPAD/5458 PAD:6055 PAD:11765 0.0375882
rPAD/5459 PAD:6055 PAD:11763 1.5
rPAD/5460 PAD:6054 PAD:6057 0.0375882
rPAD/5461 PAD:6054 PAD:6055 1.5
rPAD/5462 PAD:6052 PAD:11756 0.0375882
rPAD/5463 PAD:6052 PAD:6055 0.0751765
rPAD/5464 PAD:6052 PAD:11760 1.5
rPAD/5465 PAD:6051 PAD:6054 0.0751765
rPAD/5466 PAD:6051 PAD:6052 1.5
rPAD/5467 PAD:6048 PAD:6051 0.0375882
rPAD/5468 PAD:6048 PAD:11756 1.5
rPAD/5469 PAD:6046 PAD:11756 0.0751765
rPAD/5470 PAD:6046 PAD:11754 1.5
rPAD/5471 PAD:6045 PAD:6048 0.0751765
rPAD/5472 PAD:6045 PAD:6046 1.5
rPAD/5473 PAD:6043 PAD:6046 0.0375882
rPAD/5474 PAD:6043 PAD:11751 1.5
rPAD/5475 PAD:6042 PAD:6045 0.0375882
rPAD/5476 PAD:6042 PAD:6043 1.5
rPAD/5477 PAD:6040 PAD:6043 0.0751765
rPAD/5478 PAD:6040 PAD:11748 1.5
rPAD/5479 PAD:6039 PAD:6042 0.0751765
rPAD/5480 PAD:6039 PAD:6040 1.5
rPAD/5481 PAD:6037 PAD:6040 0.0375882
rPAD/5482 PAD:6037 PAD:11745 1.5
rPAD/5483 PAD:6036 PAD:6039 0.0375882
rPAD/5484 PAD:6036 PAD:6037 1.5
rPAD/5485 PAD:6034 PAD:6037 0.0751765
rPAD/5486 PAD:6034 PAD:11742 1.5
rPAD/5487 PAD:6033 PAD:6036 0.0751765
rPAD/5488 PAD:6033 PAD:6034 1.5
rPAD/5489 PAD:6031 PAD:11735 0.0751765
rPAD/5490 PAD:6031 PAD:6034 0.0375882
rPAD/5491 PAD:6031 PAD:11739 1.5
rPAD/5492 PAD:6030 PAD:6033 0.0375882
rPAD/5493 PAD:6030 PAD:6031 1.5
rPAD/5494 PAD:6027 PAD:6030 0.0751765
rPAD/5495 PAD:6027 PAD:11735 1.5
rPAD/5496 PAD:6025 PAD:11735 0.0375882
rPAD/5497 PAD:6025 PAD:11733 1.5
rPAD/5498 PAD:6024 PAD:6027 0.0375882
rPAD/5499 PAD:6024 PAD:6025 1.5
rPAD/5500 PAD:6022 PAD:6025 0.0751765
rPAD/5501 PAD:6022 PAD:11730 1.5
rPAD/5502 PAD:6021 PAD:6024 0.0751765
rPAD/5503 PAD:6021 PAD:6022 1.5
rPAD/5504 PAD:6019 PAD:6022 0.0375882
rPAD/5505 PAD:6019 PAD:11727 1.5
rPAD/5506 PAD:6018 PAD:6021 0.0375882
rPAD/5507 PAD:6018 PAD:6019 1.5
rPAD/5508 PAD:6016 PAD:6019 0.0751765
rPAD/5509 PAD:6016 PAD:11724 1.5
rPAD/5510 PAD:6015 PAD:6018 0.0751765
rPAD/5511 PAD:6015 PAD:6016 1.5
rPAD/5512 PAD:6013 PAD:6016 0.0375882
rPAD/5513 PAD:6013 PAD:11721 1.5
rPAD/5514 PAD:6012 PAD:6015 0.0375882
rPAD/5515 PAD:6012 PAD:6013 1.5
rPAD/5516 PAD:6010 PAD:6013 0.0751765
rPAD/5517 PAD:6010 PAD:11718 1.5
rPAD/5518 PAD:6009 PAD:6012 0.0751765
rPAD/5519 PAD:6009 PAD:6010 1.5
rPAD/5520 PAD:6007 PAD:6010 0.0375882
rPAD/5521 PAD:6007 PAD:11715 1.5
rPAD/5522 PAD:6006 PAD:6009 0.0375882
rPAD/5523 PAD:6006 PAD:6007 1.5
rPAD/5524 PAD:6004 PAD:14901 0.0283817
rPAD/5525 PAD:6004 PAD:6007 0.0751765
rPAD/5526 PAD:6004 PAD:11712 1.5
rPAD/5527 PAD:6003 PAD:9182 0.0378785
rPAD/5528 PAD:6003 PAD:6006 0.0751765
rPAD/5529 PAD:6003 PAD:6004 1.5
rPAD/5530 PAD:5999 PAD:11539 0.0100588
rPAD/5531 PAD:5999 PAD:11707 1.5
rPAD/5532 PAD:5998 PAD:9366 0.0670908
rPAD/5533 PAD:5998 PAD:5999 1.5
rPAD/5534 PAD:5996 PAD:5999 0.0751765
rPAD/5535 PAD:5996 PAD:11704 1.5
rPAD/5536 PAD:5995 PAD:5998 0.0751765
rPAD/5537 PAD:5995 PAD:5996 1.5
rPAD/5538 PAD:5993 PAD:11697 0.0751765
rPAD/5539 PAD:5993 PAD:5996 0.0375882
rPAD/5540 PAD:5993 PAD:11701 1.5
rPAD/5541 PAD:5992 PAD:5995 0.0375882
rPAD/5542 PAD:5992 PAD:5993 1.5
rPAD/5543 PAD:5989 PAD:5992 0.0751765
rPAD/5544 PAD:5989 PAD:11697 1.5
rPAD/5545 PAD:5987 PAD:11697 0.0375882
rPAD/5546 PAD:5987 PAD:11695 1.5
rPAD/5547 PAD:5986 PAD:5989 0.0375882
rPAD/5548 PAD:5986 PAD:5987 1.5
rPAD/5549 PAD:5984 PAD:5987 0.0751765
rPAD/5550 PAD:5984 PAD:11692 1.5
rPAD/5551 PAD:5983 PAD:5986 0.0751765
rPAD/5552 PAD:5983 PAD:5984 1.5
rPAD/5553 PAD:5981 PAD:5984 0.0375882
rPAD/5554 PAD:5981 PAD:11689 1.5
rPAD/5555 PAD:5980 PAD:5983 0.0375882
rPAD/5556 PAD:5980 PAD:5981 1.5
rPAD/5557 PAD:5978 PAD:5981 0.0751765
rPAD/5558 PAD:5978 PAD:11686 1.5
rPAD/5559 PAD:5977 PAD:5980 0.0751765
rPAD/5560 PAD:5977 PAD:5978 1.5
rPAD/5561 PAD:5975 PAD:5978 0.0375882
rPAD/5562 PAD:5975 PAD:11683 1.5
rPAD/5563 PAD:5974 PAD:5977 0.0375882
rPAD/5564 PAD:5974 PAD:5975 1.5
rPAD/5565 PAD:5972 PAD:5975 0.0751765
rPAD/5566 PAD:5972 PAD:11680 1.5
rPAD/5567 PAD:5971 PAD:5974 0.0751765
rPAD/5568 PAD:5971 PAD:5972 1.5
rPAD/5569 PAD:5969 PAD:5972 0.0375882
rPAD/5570 PAD:5969 PAD:11677 1.5
rPAD/5571 PAD:5968 PAD:5971 0.0375882
rPAD/5572 PAD:5968 PAD:5969 1.5
rPAD/5573 PAD:5966 PAD:5969 0.0751765
rPAD/5574 PAD:5966 PAD:11674 1.5
rPAD/5575 PAD:5965 PAD:5968 0.0751765
rPAD/5576 PAD:5965 PAD:5966 1.5
rPAD/5577 PAD:5963 PAD:5966 0.0375882
rPAD/5578 PAD:5963 PAD:11671 1.5
rPAD/5579 PAD:5962 PAD:5965 0.0375882
rPAD/5580 PAD:5962 PAD:5963 1.5
rPAD/5581 PAD:5960 PAD:5963 0.0751765
rPAD/5582 PAD:5960 PAD:11668 1.5
rPAD/5583 PAD:5959 PAD:5962 0.0751765
rPAD/5584 PAD:5959 PAD:5960 1.5
rPAD/5585 PAD:5957 PAD:11661 0.0751765
rPAD/5586 PAD:5957 PAD:5960 0.0375882
rPAD/5587 PAD:5957 PAD:11665 1.5
rPAD/5588 PAD:5956 PAD:5959 0.0375882
rPAD/5589 PAD:5956 PAD:5957 1.5
rPAD/5590 PAD:5953 PAD:5956 0.0751765
rPAD/5591 PAD:5953 PAD:11661 1.5
rPAD/5592 PAD:5951 PAD:11655 0.0751765
rPAD/5593 PAD:5951 PAD:11661 0.0375882
rPAD/5594 PAD:5951 PAD:11659 1.5
rPAD/5595 PAD:5950 PAD:5953 0.0375882
rPAD/5596 PAD:5950 PAD:5951 1.5
rPAD/5597 PAD:5947 PAD:5950 0.0751765
rPAD/5598 PAD:5947 PAD:11655 1.5
rPAD/5599 PAD:5944 PAD:5947 0.0375882
rPAD/5600 PAD:5944 PAD:11652 1.5
rPAD/5601 PAD:5941 PAD:5944 0.0751765
rPAD/5602 PAD:5941 PAD:11649 1.5
rPAD/5603 PAD:5939 PAD:11643 0.0751765
rPAD/5604 PAD:5939 PAD:11649 0.0375882
rPAD/5605 PAD:5939 PAD:11647 1.5
rPAD/5606 PAD:5938 PAD:5941 0.0375882
rPAD/5607 PAD:5938 PAD:5939 1.5
rPAD/5608 PAD:5935 PAD:5938 0.0751765
rPAD/5609 PAD:5935 PAD:11643 1.5
rPAD/5610 PAD:5932 PAD:5935 0.0375882
rPAD/5611 PAD:5932 PAD:11640 1.5
rPAD/5612 PAD:5930 PAD:11640 0.0751765
rPAD/5613 PAD:5930 PAD:11638 1.5
rPAD/5614 PAD:5929 PAD:5932 0.0751765
rPAD/5615 PAD:5929 PAD:5930 1.5
rPAD/5616 PAD:5927 PAD:5930 0.0375882
rPAD/5617 PAD:5927 PAD:11635 1.5
rPAD/5618 PAD:5926 PAD:5929 0.0375882
rPAD/5619 PAD:5926 PAD:5927 1.5
rPAD/5620 PAD:5924 PAD:5927 0.0751765
rPAD/5621 PAD:5924 PAD:11632 1.5
rPAD/5622 PAD:5923 PAD:5926 0.0751765
rPAD/5623 PAD:5923 PAD:5924 1.5
rPAD/5624 PAD:5921 PAD:5924 0.0375882
rPAD/5625 PAD:5921 PAD:11629 1.5
rPAD/5626 PAD:5920 PAD:5923 0.0375882
rPAD/5627 PAD:5920 PAD:5921 1.5
rPAD/5628 PAD:5918 PAD:5921 0.0751765
rPAD/5629 PAD:5918 PAD:11626 1.5
rPAD/5630 PAD:5917 PAD:5920 0.0751765
rPAD/5631 PAD:5917 PAD:5918 1.5
rPAD/5632 PAD:5915 PAD:11619 0.0751765
rPAD/5633 PAD:5915 PAD:5918 0.0375882
rPAD/5634 PAD:5915 PAD:11623 1.5
rPAD/5635 PAD:5914 PAD:5917 0.0375882
rPAD/5636 PAD:5914 PAD:5915 1.5
rPAD/5637 PAD:5911 PAD:5914 0.0751765
rPAD/5638 PAD:5911 PAD:11619 1.5
rPAD/5639 PAD:5909 PAD:11619 0.0375882
rPAD/5640 PAD:5909 PAD:11617 1.5
rPAD/5641 PAD:5908 PAD:5911 0.0375882
rPAD/5642 PAD:5908 PAD:5909 1.5
rPAD/5643 PAD:5906 PAD:5909 0.0751765
rPAD/5644 PAD:5906 PAD:11614 1.5
rPAD/5645 PAD:5905 PAD:5908 0.0751765
rPAD/5646 PAD:5905 PAD:5906 1.5
rPAD/5647 PAD:5903 PAD:11607 0.0751765
rPAD/5648 PAD:5903 PAD:5906 0.0375882
rPAD/5649 PAD:5903 PAD:11611 1.5
rPAD/5650 PAD:5902 PAD:5905 0.0375882
rPAD/5651 PAD:5902 PAD:5903 1.5
rPAD/5652 PAD:5899 PAD:5902 0.0751765
rPAD/5653 PAD:5899 PAD:11607 1.5
rPAD/5654 PAD:5896 PAD:5899 0.0375882
rPAD/5655 PAD:5896 PAD:11604 1.5
rPAD/5656 PAD:5893 PAD:5896 0.0751765
rPAD/5657 PAD:5893 PAD:11601 1.5
rPAD/5658 PAD:5890 PAD:5893 0.0375882
rPAD/5659 PAD:5890 PAD:11598 1.5
rPAD/5660 PAD:5887 PAD:5890 0.0751765
rPAD/5661 PAD:5887 PAD:11595 1.5
rPAD/5662 PAD:5885 PAD:11595 0.0375882
rPAD/5663 PAD:5885 PAD:11593 1.5
rPAD/5664 PAD:5884 PAD:5887 0.0375882
rPAD/5665 PAD:5884 PAD:5885 1.5
rPAD/5666 PAD:5882 PAD:11586 0.0375882
rPAD/5667 PAD:5882 PAD:5885 0.0751765
rPAD/5668 PAD:5882 PAD:11590 1.5
rPAD/5669 PAD:5881 PAD:5884 0.0751765
rPAD/5670 PAD:5881 PAD:5882 1.5
rPAD/5671 PAD:5878 PAD:5881 0.0375882
rPAD/5672 PAD:5878 PAD:11586 1.5
rPAD/5673 PAD:5876 PAD:11586 0.0751765
rPAD/5674 PAD:5876 PAD:11584 1.5
rPAD/5675 PAD:5875 PAD:5878 0.0751765
rPAD/5676 PAD:5875 PAD:5876 1.5
rPAD/5677 PAD:5873 PAD:5876 0.0375882
rPAD/5678 PAD:5873 PAD:11581 1.5
rPAD/5679 PAD:5872 PAD:5875 0.0375882
rPAD/5680 PAD:5872 PAD:5873 1.5
rPAD/5681 PAD:5870 PAD:5873 0.0751765
rPAD/5682 PAD:5870 PAD:11578 1.5
rPAD/5683 PAD:5869 PAD:5872 0.0751765
rPAD/5684 PAD:5869 PAD:5870 1.5
rPAD/5685 PAD:5867 PAD:5870 0.0375882
rPAD/5686 PAD:5867 PAD:11575 1.5
rPAD/5687 PAD:5866 PAD:5869 0.0375882
rPAD/5688 PAD:5866 PAD:5867 1.5
rPAD/5689 PAD:5864 PAD:5867 0.0751765
rPAD/5690 PAD:5864 PAD:11572 1.5
rPAD/5691 PAD:5863 PAD:5866 0.0751765
rPAD/5692 PAD:5863 PAD:5864 1.5
rPAD/5693 PAD:5861 PAD:11565 0.0751765
rPAD/5694 PAD:5861 PAD:5864 0.0375882
rPAD/5695 PAD:5861 PAD:11569 1.5
rPAD/5696 PAD:5860 PAD:5863 0.0375882
rPAD/5697 PAD:5860 PAD:5861 1.5
rPAD/5698 PAD:5857 PAD:5860 0.0751765
rPAD/5699 PAD:5857 PAD:11565 1.5
rPAD/5700 PAD:5855 PAD:11565 0.0375882
rPAD/5701 PAD:5855 PAD:11563 1.5
rPAD/5702 PAD:5854 PAD:5857 0.0375882
rPAD/5703 PAD:5854 PAD:5855 1.5
rPAD/5704 PAD:5852 PAD:5855 0.0751765
rPAD/5705 PAD:5852 PAD:11560 1.5
rPAD/5706 PAD:5851 PAD:5854 0.0751765
rPAD/5707 PAD:5851 PAD:5852 1.5
rPAD/5708 PAD:5849 PAD:5852 0.0375882
rPAD/5709 PAD:5849 PAD:11557 1.5
rPAD/5710 PAD:5848 PAD:5851 0.0375882
rPAD/5711 PAD:5848 PAD:5849 1.5
rPAD/5712 PAD:5846 PAD:5849 0.0751765
rPAD/5713 PAD:5846 PAD:11554 1.5
rPAD/5714 PAD:5845 PAD:5848 0.0751765
rPAD/5715 PAD:5845 PAD:5846 1.5
rPAD/5716 PAD:5843 PAD:5846 0.0375882
rPAD/5717 PAD:5843 PAD:11551 1.5
rPAD/5718 PAD:5842 PAD:5845 0.0375882
rPAD/5719 PAD:5842 PAD:5843 1.5
rPAD/5720 PAD:5840 PAD:5843 0.0751765
rPAD/5721 PAD:5840 PAD:11548 1.5
rPAD/5722 PAD:5839 PAD:5842 0.0751765
rPAD/5723 PAD:5839 PAD:5840 1.5
rPAD/5724 PAD:5837 PAD:5840 0.0375882
rPAD/5725 PAD:5837 PAD:11545 1.5
rPAD/5726 PAD:5836 PAD:5839 0.0375882
rPAD/5727 PAD:5836 PAD:5837 1.5
rPAD/5728 PAD:5834 PAD:14895 0.0283817
rPAD/5729 PAD:5834 PAD:5837 0.0751765
rPAD/5730 PAD:5834 PAD:11542 1.5
rPAD/5731 PAD:5833 PAD:9175 0.0378785
rPAD/5732 PAD:5833 PAD:5836 0.0751765
rPAD/5733 PAD:5833 PAD:5834 1.5
rPAD/5734 PAD:5829 PAD:11369 0.0100588
rPAD/5735 PAD:5829 PAD:11537 1.5
rPAD/5736 PAD:5828 PAD:9362 0.0670908
rPAD/5737 PAD:5828 PAD:5829 1.5
rPAD/5738 PAD:5826 PAD:5829 0.0751765
rPAD/5739 PAD:5826 PAD:11534 1.5
rPAD/5740 PAD:5825 PAD:5828 0.0751765
rPAD/5741 PAD:5825 PAD:5826 1.5
rPAD/5742 PAD:5823 PAD:11527 0.0751765
rPAD/5743 PAD:5823 PAD:5826 0.0375882
rPAD/5744 PAD:5823 PAD:11531 1.5
rPAD/5745 PAD:5822 PAD:5825 0.0375882
rPAD/5746 PAD:5822 PAD:5823 1.5
rPAD/5747 PAD:5819 PAD:5822 0.0751765
rPAD/5748 PAD:5819 PAD:11527 1.5
rPAD/5749 PAD:5817 PAD:11527 0.0375882
rPAD/5750 PAD:5817 PAD:11525 1.5
rPAD/5751 PAD:5816 PAD:5819 0.0375882
rPAD/5752 PAD:5816 PAD:5817 1.5
rPAD/5753 PAD:5814 PAD:5817 0.0751765
rPAD/5754 PAD:5814 PAD:11522 1.5
rPAD/5755 PAD:5813 PAD:5816 0.0751765
rPAD/5756 PAD:5813 PAD:5814 1.5
rPAD/5757 PAD:5811 PAD:5814 0.0375882
rPAD/5758 PAD:5811 PAD:11519 1.5
rPAD/5759 PAD:5810 PAD:5813 0.0375882
rPAD/5760 PAD:5810 PAD:5811 1.5
rPAD/5761 PAD:5808 PAD:5811 0.0751765
rPAD/5762 PAD:5808 PAD:11516 1.5
rPAD/5763 PAD:5807 PAD:5810 0.0751765
rPAD/5764 PAD:5807 PAD:5808 1.5
rPAD/5765 PAD:5805 PAD:5808 0.0375882
rPAD/5766 PAD:5805 PAD:11513 1.5
rPAD/5767 PAD:5804 PAD:5807 0.0375882
rPAD/5768 PAD:5804 PAD:5805 1.5
rPAD/5769 PAD:5802 PAD:5805 0.0751765
rPAD/5770 PAD:5802 PAD:11510 1.5
rPAD/5771 PAD:5801 PAD:5804 0.0751765
rPAD/5772 PAD:5801 PAD:5802 1.5
rPAD/5773 PAD:5799 PAD:5802 0.0375882
rPAD/5774 PAD:5799 PAD:11507 1.5
rPAD/5775 PAD:5798 PAD:5801 0.0375882
rPAD/5776 PAD:5798 PAD:5799 1.5
rPAD/5777 PAD:5796 PAD:5799 0.0751765
rPAD/5778 PAD:5796 PAD:11504 1.5
rPAD/5779 PAD:5795 PAD:5798 0.0751765
rPAD/5780 PAD:5795 PAD:5796 1.5
rPAD/5781 PAD:5793 PAD:5796 0.0375882
rPAD/5782 PAD:5793 PAD:11501 1.5
rPAD/5783 PAD:5792 PAD:5795 0.0375882
rPAD/5784 PAD:5792 PAD:5793 1.5
rPAD/5785 PAD:5790 PAD:5793 0.0751765
rPAD/5786 PAD:5790 PAD:11498 1.5
rPAD/5787 PAD:5789 PAD:5792 0.0751765
rPAD/5788 PAD:5789 PAD:5790 1.5
rPAD/5789 PAD:5787 PAD:11491 0.0751765
rPAD/5790 PAD:5787 PAD:5790 0.0375882
rPAD/5791 PAD:5787 PAD:11495 1.5
rPAD/5792 PAD:5786 PAD:5789 0.0375882
rPAD/5793 PAD:5786 PAD:5787 1.5
rPAD/5794 PAD:5783 PAD:5786 0.0751765
rPAD/5795 PAD:5783 PAD:11491 1.5
rPAD/5796 PAD:5781 PAD:11485 0.0751765
rPAD/5797 PAD:5781 PAD:11491 0.0375882
rPAD/5798 PAD:5781 PAD:11489 1.5
rPAD/5799 PAD:5780 PAD:5783 0.0375882
rPAD/5800 PAD:5780 PAD:5781 1.5
rPAD/5801 PAD:5777 PAD:5780 0.0751765
rPAD/5802 PAD:5777 PAD:11485 1.5
rPAD/5803 PAD:5774 PAD:5777 0.0375882
rPAD/5804 PAD:5774 PAD:11482 1.5
rPAD/5805 PAD:5771 PAD:5774 0.0751765
rPAD/5806 PAD:5771 PAD:11479 1.5
rPAD/5807 PAD:5769 PAD:11473 0.0751765
rPAD/5808 PAD:5769 PAD:11479 0.0375882
rPAD/5809 PAD:5769 PAD:11477 1.5
rPAD/5810 PAD:5768 PAD:5771 0.0375882
rPAD/5811 PAD:5768 PAD:5769 1.5
rPAD/5812 PAD:5765 PAD:5768 0.0751765
rPAD/5813 PAD:5765 PAD:11473 1.5
rPAD/5814 PAD:5762 PAD:5765 0.0375882
rPAD/5815 PAD:5762 PAD:11470 1.5
rPAD/5816 PAD:5760 PAD:11470 0.0751765
rPAD/5817 PAD:5760 PAD:11468 1.5
rPAD/5818 PAD:5759 PAD:5762 0.0751765
rPAD/5819 PAD:5759 PAD:5760 1.5
rPAD/5820 PAD:5757 PAD:5760 0.0375882
rPAD/5821 PAD:5757 PAD:11465 1.5
rPAD/5822 PAD:5756 PAD:5759 0.0375882
rPAD/5823 PAD:5756 PAD:5757 1.5
rPAD/5824 PAD:5754 PAD:5757 0.0751765
rPAD/5825 PAD:5754 PAD:11462 1.5
rPAD/5826 PAD:5753 PAD:5756 0.0751765
rPAD/5827 PAD:5753 PAD:5754 1.5
rPAD/5828 PAD:5751 PAD:5754 0.0375882
rPAD/5829 PAD:5751 PAD:11459 1.5
rPAD/5830 PAD:5750 PAD:5753 0.0375882
rPAD/5831 PAD:5750 PAD:5751 1.5
rPAD/5832 PAD:5748 PAD:5751 0.0751765
rPAD/5833 PAD:5748 PAD:11456 1.5
rPAD/5834 PAD:5747 PAD:5750 0.0751765
rPAD/5835 PAD:5747 PAD:5748 1.5
rPAD/5836 PAD:5745 PAD:11449 0.0751765
rPAD/5837 PAD:5745 PAD:5748 0.0375882
rPAD/5838 PAD:5745 PAD:11453 1.5
rPAD/5839 PAD:5744 PAD:5747 0.0375882
rPAD/5840 PAD:5744 PAD:5745 1.5
rPAD/5841 PAD:5741 PAD:5744 0.0751765
rPAD/5842 PAD:5741 PAD:11449 1.5
rPAD/5843 PAD:5739 PAD:11449 0.0375882
rPAD/5844 PAD:5739 PAD:11447 1.5
rPAD/5845 PAD:5738 PAD:5741 0.0375882
rPAD/5846 PAD:5738 PAD:5739 1.5
rPAD/5847 PAD:5736 PAD:5739 0.0751765
rPAD/5848 PAD:5736 PAD:11444 1.5
rPAD/5849 PAD:5735 PAD:5738 0.0751765
rPAD/5850 PAD:5735 PAD:5736 1.5
rPAD/5851 PAD:5733 PAD:11437 0.0751765
rPAD/5852 PAD:5733 PAD:5736 0.0375882
rPAD/5853 PAD:5733 PAD:11441 1.5
rPAD/5854 PAD:5732 PAD:5735 0.0375882
rPAD/5855 PAD:5732 PAD:5733 1.5
rPAD/5856 PAD:5729 PAD:5732 0.0751765
rPAD/5857 PAD:5729 PAD:11437 1.5
rPAD/5858 PAD:5726 PAD:5729 0.0375882
rPAD/5859 PAD:5726 PAD:11434 1.5
rPAD/5860 PAD:5723 PAD:5726 0.0751765
rPAD/5861 PAD:5723 PAD:11431 1.5
rPAD/5862 PAD:5720 PAD:5723 0.0375882
rPAD/5863 PAD:5720 PAD:11428 1.5
rPAD/5864 PAD:5717 PAD:5720 0.0751765
rPAD/5865 PAD:5717 PAD:11425 1.5
rPAD/5866 PAD:5715 PAD:11425 0.0375882
rPAD/5867 PAD:5715 PAD:11423 1.5
rPAD/5868 PAD:5714 PAD:5717 0.0375882
rPAD/5869 PAD:5714 PAD:5715 1.5
rPAD/5870 PAD:5712 PAD:11416 0.0375882
rPAD/5871 PAD:5712 PAD:5715 0.0751765
rPAD/5872 PAD:5712 PAD:11420 1.5
rPAD/5873 PAD:5711 PAD:5714 0.0751765
rPAD/5874 PAD:5711 PAD:5712 1.5
rPAD/5875 PAD:5708 PAD:5711 0.0375882
rPAD/5876 PAD:5708 PAD:11416 1.5
rPAD/5877 PAD:5706 PAD:11416 0.0751765
rPAD/5878 PAD:5706 PAD:11414 1.5
rPAD/5879 PAD:5705 PAD:5708 0.0751765
rPAD/5880 PAD:5705 PAD:5706 1.5
rPAD/5881 PAD:5703 PAD:5706 0.0375882
rPAD/5882 PAD:5703 PAD:11411 1.5
rPAD/5883 PAD:5702 PAD:5705 0.0375882
rPAD/5884 PAD:5702 PAD:5703 1.5
rPAD/5885 PAD:5700 PAD:5703 0.0751765
rPAD/5886 PAD:5700 PAD:11408 1.5
rPAD/5887 PAD:5699 PAD:5702 0.0751765
rPAD/5888 PAD:5699 PAD:5700 1.5
rPAD/5889 PAD:5697 PAD:5700 0.0375882
rPAD/5890 PAD:5697 PAD:11405 1.5
rPAD/5891 PAD:5696 PAD:5699 0.0375882
rPAD/5892 PAD:5696 PAD:5697 1.5
rPAD/5893 PAD:5694 PAD:5697 0.0751765
rPAD/5894 PAD:5694 PAD:11402 1.5
rPAD/5895 PAD:5693 PAD:5696 0.0751765
rPAD/5896 PAD:5693 PAD:5694 1.5
rPAD/5897 PAD:5691 PAD:11395 0.0751765
rPAD/5898 PAD:5691 PAD:5694 0.0375882
rPAD/5899 PAD:5691 PAD:11399 1.5
rPAD/5900 PAD:5690 PAD:5693 0.0375882
rPAD/5901 PAD:5690 PAD:5691 1.5
rPAD/5902 PAD:5687 PAD:5690 0.0751765
rPAD/5903 PAD:5687 PAD:11395 1.5
rPAD/5904 PAD:5685 PAD:11395 0.0375882
rPAD/5905 PAD:5685 PAD:11393 1.5
rPAD/5906 PAD:5684 PAD:5687 0.0375882
rPAD/5907 PAD:5684 PAD:5685 1.5
rPAD/5908 PAD:5682 PAD:5685 0.0751765
rPAD/5909 PAD:5682 PAD:11390 1.5
rPAD/5910 PAD:5681 PAD:5684 0.0751765
rPAD/5911 PAD:5681 PAD:5682 1.5
rPAD/5912 PAD:5679 PAD:5682 0.0375882
rPAD/5913 PAD:5679 PAD:11387 1.5
rPAD/5914 PAD:5678 PAD:5681 0.0375882
rPAD/5915 PAD:5678 PAD:5679 1.5
rPAD/5916 PAD:5676 PAD:5679 0.0751765
rPAD/5917 PAD:5676 PAD:11384 1.5
rPAD/5918 PAD:5675 PAD:5678 0.0751765
rPAD/5919 PAD:5675 PAD:5676 1.5
rPAD/5920 PAD:5673 PAD:5676 0.0375882
rPAD/5921 PAD:5673 PAD:11381 1.5
rPAD/5922 PAD:5672 PAD:5675 0.0375882
rPAD/5923 PAD:5672 PAD:5673 1.5
rPAD/5924 PAD:5670 PAD:5673 0.0751765
rPAD/5925 PAD:5670 PAD:11378 1.5
rPAD/5926 PAD:5669 PAD:5672 0.0751765
rPAD/5927 PAD:5669 PAD:5670 1.5
rPAD/5928 PAD:5667 PAD:5670 0.0375882
rPAD/5929 PAD:5667 PAD:11375 1.5
rPAD/5930 PAD:5666 PAD:5669 0.0375882
rPAD/5931 PAD:5666 PAD:5667 1.5
rPAD/5932 PAD:5664 PAD:14887 0.0283817
rPAD/5933 PAD:5664 PAD:5667 0.0751765
rPAD/5934 PAD:5664 PAD:11372 1.5
rPAD/5935 PAD:5663 PAD:9168 0.0378785
rPAD/5936 PAD:5663 PAD:5666 0.0751765
rPAD/5937 PAD:5663 PAD:5664 1.5
rPAD/5938 PAD:5659 PAD:11199 0.0100588
rPAD/5939 PAD:5659 PAD:11367 1.5
rPAD/5940 PAD:5658 PAD:9357 0.0670908
rPAD/5941 PAD:5658 PAD:5659 1.5
rPAD/5942 PAD:5656 PAD:5659 0.0751765
rPAD/5943 PAD:5656 PAD:11364 1.5
rPAD/5944 PAD:5655 PAD:5658 0.0751765
rPAD/5945 PAD:5655 PAD:5656 1.5
rPAD/5946 PAD:5653 PAD:11357 0.0751765
rPAD/5947 PAD:5653 PAD:5656 0.0375882
rPAD/5948 PAD:5653 PAD:11361 1.5
rPAD/5949 PAD:5652 PAD:5655 0.0375882
rPAD/5950 PAD:5652 PAD:5653 1.5
rPAD/5951 PAD:5649 PAD:5652 0.0751765
rPAD/5952 PAD:5649 PAD:11357 1.5
rPAD/5953 PAD:5647 PAD:11357 0.0375882
rPAD/5954 PAD:5647 PAD:11355 1.5
rPAD/5955 PAD:5646 PAD:5649 0.0375882
rPAD/5956 PAD:5646 PAD:5647 1.5
rPAD/5957 PAD:5644 PAD:5647 0.0751765
rPAD/5958 PAD:5644 PAD:11352 1.5
rPAD/5959 PAD:5643 PAD:5646 0.0751765
rPAD/5960 PAD:5643 PAD:5644 1.5
rPAD/5961 PAD:5641 PAD:5644 0.0375882
rPAD/5962 PAD:5641 PAD:11349 1.5
rPAD/5963 PAD:5640 PAD:5643 0.0375882
rPAD/5964 PAD:5640 PAD:5641 1.5
rPAD/5965 PAD:5638 PAD:5641 0.0751765
rPAD/5966 PAD:5638 PAD:11346 1.5
rPAD/5967 PAD:5637 PAD:5640 0.0751765
rPAD/5968 PAD:5637 PAD:5638 1.5
rPAD/5969 PAD:5635 PAD:5638 0.0375882
rPAD/5970 PAD:5635 PAD:11343 1.5
rPAD/5971 PAD:5634 PAD:5637 0.0375882
rPAD/5972 PAD:5634 PAD:5635 1.5
rPAD/5973 PAD:5632 PAD:5635 0.0751765
rPAD/5974 PAD:5632 PAD:11340 1.5
rPAD/5975 PAD:5631 PAD:5634 0.0751765
rPAD/5976 PAD:5631 PAD:5632 1.5
rPAD/5977 PAD:5629 PAD:5632 0.0375882
rPAD/5978 PAD:5629 PAD:11337 1.5
rPAD/5979 PAD:5628 PAD:5631 0.0375882
rPAD/5980 PAD:5628 PAD:5629 1.5
rPAD/5981 PAD:5626 PAD:5629 0.0751765
rPAD/5982 PAD:5626 PAD:11334 1.5
rPAD/5983 PAD:5625 PAD:5628 0.0751765
rPAD/5984 PAD:5625 PAD:5626 1.5
rPAD/5985 PAD:5623 PAD:5626 0.0375882
rPAD/5986 PAD:5623 PAD:11331 1.5
rPAD/5987 PAD:5622 PAD:5625 0.0375882
rPAD/5988 PAD:5622 PAD:5623 1.5
rPAD/5989 PAD:5620 PAD:5623 0.0751765
rPAD/5990 PAD:5620 PAD:11328 1.5
rPAD/5991 PAD:5619 PAD:5622 0.0751765
rPAD/5992 PAD:5619 PAD:5620 1.5
rPAD/5993 PAD:5617 PAD:11321 0.0751765
rPAD/5994 PAD:5617 PAD:5620 0.0375882
rPAD/5995 PAD:5617 PAD:11325 1.5
rPAD/5996 PAD:5616 PAD:5619 0.0375882
rPAD/5997 PAD:5616 PAD:5617 1.5
rPAD/5998 PAD:5613 PAD:5616 0.0751765
rPAD/5999 PAD:5613 PAD:11321 1.5
rPAD/6000 PAD:5611 PAD:11315 0.0751765
rPAD/6001 PAD:5611 PAD:11321 0.0375882
rPAD/6002 PAD:5611 PAD:11319 1.5
rPAD/6003 PAD:5610 PAD:5613 0.0375882
rPAD/6004 PAD:5610 PAD:5611 1.5
rPAD/6005 PAD:5607 PAD:5610 0.0751765
rPAD/6006 PAD:5607 PAD:11315 1.5
rPAD/6007 PAD:5604 PAD:5607 0.0375882
rPAD/6008 PAD:5604 PAD:11312 1.5
rPAD/6009 PAD:5601 PAD:5604 0.0751765
rPAD/6010 PAD:5601 PAD:11309 1.5
rPAD/6011 PAD:5599 PAD:11303 0.0751765
rPAD/6012 PAD:5599 PAD:11309 0.0375882
rPAD/6013 PAD:5599 PAD:11307 1.5
rPAD/6014 PAD:5598 PAD:5601 0.0375882
rPAD/6015 PAD:5598 PAD:5599 1.5
rPAD/6016 PAD:5595 PAD:5598 0.0751765
rPAD/6017 PAD:5595 PAD:11303 1.5
rPAD/6018 PAD:5592 PAD:5595 0.0375882
rPAD/6019 PAD:5592 PAD:11300 1.5
rPAD/6020 PAD:5590 PAD:11300 0.0751765
rPAD/6021 PAD:5590 PAD:11298 1.5
rPAD/6022 PAD:5589 PAD:5592 0.0751765
rPAD/6023 PAD:5589 PAD:5590 1.5
rPAD/6024 PAD:5587 PAD:5590 0.0375882
rPAD/6025 PAD:5587 PAD:11295 1.5
rPAD/6026 PAD:5586 PAD:5589 0.0375882
rPAD/6027 PAD:5586 PAD:5587 1.5
rPAD/6028 PAD:5584 PAD:5587 0.0751765
rPAD/6029 PAD:5584 PAD:11292 1.5
rPAD/6030 PAD:5583 PAD:5586 0.0751765
rPAD/6031 PAD:5583 PAD:5584 1.5
rPAD/6032 PAD:5581 PAD:5584 0.0375882
rPAD/6033 PAD:5581 PAD:11289 1.5
rPAD/6034 PAD:5580 PAD:5583 0.0375882
rPAD/6035 PAD:5580 PAD:5581 1.5
rPAD/6036 PAD:5578 PAD:5581 0.0751765
rPAD/6037 PAD:5578 PAD:11286 1.5
rPAD/6038 PAD:5577 PAD:5580 0.0751765
rPAD/6039 PAD:5577 PAD:5578 1.5
rPAD/6040 PAD:5575 PAD:11279 0.0751765
rPAD/6041 PAD:5575 PAD:5578 0.0375882
rPAD/6042 PAD:5575 PAD:11283 1.5
rPAD/6043 PAD:5574 PAD:5577 0.0375882
rPAD/6044 PAD:5574 PAD:5575 1.5
rPAD/6045 PAD:5571 PAD:5574 0.0751765
rPAD/6046 PAD:5571 PAD:11279 1.5
rPAD/6047 PAD:5569 PAD:11279 0.0375882
rPAD/6048 PAD:5569 PAD:11277 1.5
rPAD/6049 PAD:5568 PAD:5571 0.0375882
rPAD/6050 PAD:5568 PAD:5569 1.5
rPAD/6051 PAD:5566 PAD:5569 0.0751765
rPAD/6052 PAD:5566 PAD:11274 1.5
rPAD/6053 PAD:5565 PAD:5568 0.0751765
rPAD/6054 PAD:5565 PAD:5566 1.5
rPAD/6055 PAD:5563 PAD:11267 0.0751765
rPAD/6056 PAD:5563 PAD:5566 0.0375882
rPAD/6057 PAD:5563 PAD:11271 1.5
rPAD/6058 PAD:5562 PAD:5565 0.0375882
rPAD/6059 PAD:5562 PAD:5563 1.5
rPAD/6060 PAD:5559 PAD:5562 0.0751765
rPAD/6061 PAD:5559 PAD:11267 1.5
rPAD/6062 PAD:5556 PAD:5559 0.0375882
rPAD/6063 PAD:5556 PAD:11264 1.5
rPAD/6064 PAD:5553 PAD:5556 0.0751765
rPAD/6065 PAD:5553 PAD:11261 1.5
rPAD/6066 PAD:5550 PAD:5553 0.0375882
rPAD/6067 PAD:5550 PAD:11258 1.5
rPAD/6068 PAD:5547 PAD:5550 0.0751765
rPAD/6069 PAD:5547 PAD:11255 1.5
rPAD/6070 PAD:5545 PAD:11255 0.0375882
rPAD/6071 PAD:5545 PAD:11253 1.5
rPAD/6072 PAD:5544 PAD:5547 0.0375882
rPAD/6073 PAD:5544 PAD:5545 1.5
rPAD/6074 PAD:5542 PAD:11246 0.0375882
rPAD/6075 PAD:5542 PAD:5545 0.0751765
rPAD/6076 PAD:5542 PAD:11250 1.5
rPAD/6077 PAD:5541 PAD:5544 0.0751765
rPAD/6078 PAD:5541 PAD:5542 1.5
rPAD/6079 PAD:5538 PAD:5541 0.0375882
rPAD/6080 PAD:5538 PAD:11246 1.5
rPAD/6081 PAD:5536 PAD:11246 0.0751765
rPAD/6082 PAD:5536 PAD:11244 1.5
rPAD/6083 PAD:5535 PAD:5538 0.0751765
rPAD/6084 PAD:5535 PAD:5536 1.5
rPAD/6085 PAD:5533 PAD:5536 0.0375882
rPAD/6086 PAD:5533 PAD:11241 1.5
rPAD/6087 PAD:5532 PAD:5535 0.0375882
rPAD/6088 PAD:5532 PAD:5533 1.5
rPAD/6089 PAD:5530 PAD:5533 0.0751765
rPAD/6090 PAD:5530 PAD:11238 1.5
rPAD/6091 PAD:5529 PAD:5532 0.0751765
rPAD/6092 PAD:5529 PAD:5530 1.5
rPAD/6093 PAD:5527 PAD:5530 0.0375882
rPAD/6094 PAD:5527 PAD:11235 1.5
rPAD/6095 PAD:5526 PAD:5529 0.0375882
rPAD/6096 PAD:5526 PAD:5527 1.5
rPAD/6097 PAD:5524 PAD:5527 0.0751765
rPAD/6098 PAD:5524 PAD:11232 1.5
rPAD/6099 PAD:5523 PAD:5526 0.0751765
rPAD/6100 PAD:5523 PAD:5524 1.5
rPAD/6101 PAD:5521 PAD:11225 0.0751765
rPAD/6102 PAD:5521 PAD:5524 0.0375882
rPAD/6103 PAD:5521 PAD:11229 1.5
rPAD/6104 PAD:5520 PAD:5523 0.0375882
rPAD/6105 PAD:5520 PAD:5521 1.5
rPAD/6106 PAD:5517 PAD:5520 0.0751765
rPAD/6107 PAD:5517 PAD:11225 1.5
rPAD/6108 PAD:5515 PAD:11225 0.0375882
rPAD/6109 PAD:5515 PAD:11223 1.5
rPAD/6110 PAD:5514 PAD:5517 0.0375882
rPAD/6111 PAD:5514 PAD:5515 1.5
rPAD/6112 PAD:5512 PAD:5515 0.0751765
rPAD/6113 PAD:5512 PAD:11220 1.5
rPAD/6114 PAD:5511 PAD:5514 0.0751765
rPAD/6115 PAD:5511 PAD:5512 1.5
rPAD/6116 PAD:5509 PAD:5512 0.0375882
rPAD/6117 PAD:5509 PAD:11217 1.5
rPAD/6118 PAD:5508 PAD:5511 0.0375882
rPAD/6119 PAD:5508 PAD:5509 1.5
rPAD/6120 PAD:5506 PAD:5509 0.0751765
rPAD/6121 PAD:5506 PAD:11214 1.5
rPAD/6122 PAD:5505 PAD:5508 0.0751765
rPAD/6123 PAD:5505 PAD:5506 1.5
rPAD/6124 PAD:5503 PAD:5506 0.0375882
rPAD/6125 PAD:5503 PAD:11211 1.5
rPAD/6126 PAD:5502 PAD:5505 0.0375882
rPAD/6127 PAD:5502 PAD:5503 1.5
rPAD/6128 PAD:5500 PAD:5503 0.0751765
rPAD/6129 PAD:5500 PAD:11208 1.5
rPAD/6130 PAD:5499 PAD:5502 0.0751765
rPAD/6131 PAD:5499 PAD:5500 1.5
rPAD/6132 PAD:5497 PAD:5500 0.0375882
rPAD/6133 PAD:5497 PAD:11205 1.5
rPAD/6134 PAD:5496 PAD:5499 0.0375882
rPAD/6135 PAD:5496 PAD:5497 1.5
rPAD/6136 PAD:5494 PAD:14885 0.0283817
rPAD/6137 PAD:5494 PAD:5497 0.0751765
rPAD/6138 PAD:5494 PAD:11202 1.5
rPAD/6139 PAD:5493 PAD:9164 0.0378785
rPAD/6140 PAD:5493 PAD:5496 0.0751765
rPAD/6141 PAD:5493 PAD:5494 1.5
rPAD/6142 PAD:5489 PAD:11029 0.0100588
rPAD/6143 PAD:5489 PAD:11197 1.5
rPAD/6144 PAD:5488 PAD:9353 0.0670908
rPAD/6145 PAD:5488 PAD:5489 1.5
rPAD/6146 PAD:5486 PAD:5489 0.0751765
rPAD/6147 PAD:5486 PAD:11194 1.5
rPAD/6148 PAD:5485 PAD:5488 0.0751765
rPAD/6149 PAD:5485 PAD:5486 1.5
rPAD/6150 PAD:5483 PAD:11187 0.0751765
rPAD/6151 PAD:5483 PAD:5486 0.0375882
rPAD/6152 PAD:5483 PAD:11191 1.5
rPAD/6153 PAD:5482 PAD:5485 0.0375882
rPAD/6154 PAD:5482 PAD:5483 1.5
rPAD/6155 PAD:5479 PAD:5482 0.0751765
rPAD/6156 PAD:5479 PAD:11187 1.5
rPAD/6157 PAD:5477 PAD:11187 0.0375882
rPAD/6158 PAD:5477 PAD:11185 1.5
rPAD/6159 PAD:5476 PAD:5479 0.0375882
rPAD/6160 PAD:5476 PAD:5477 1.5
rPAD/6161 PAD:5474 PAD:5477 0.0751765
rPAD/6162 PAD:5474 PAD:11182 1.5
rPAD/6163 PAD:5473 PAD:5476 0.0751765
rPAD/6164 PAD:5473 PAD:5474 1.5
rPAD/6165 PAD:5471 PAD:5474 0.0375882
rPAD/6166 PAD:5471 PAD:11179 1.5
rPAD/6167 PAD:5470 PAD:5473 0.0375882
rPAD/6168 PAD:5470 PAD:5471 1.5
rPAD/6169 PAD:5468 PAD:5471 0.0751765
rPAD/6170 PAD:5468 PAD:11176 1.5
rPAD/6171 PAD:5467 PAD:5470 0.0751765
rPAD/6172 PAD:5467 PAD:5468 1.5
rPAD/6173 PAD:5465 PAD:5468 0.0375882
rPAD/6174 PAD:5465 PAD:11173 1.5
rPAD/6175 PAD:5464 PAD:5467 0.0375882
rPAD/6176 PAD:5464 PAD:5465 1.5
rPAD/6177 PAD:5462 PAD:5465 0.0751765
rPAD/6178 PAD:5462 PAD:11170 1.5
rPAD/6179 PAD:5461 PAD:5464 0.0751765
rPAD/6180 PAD:5461 PAD:5462 1.5
rPAD/6181 PAD:5459 PAD:5462 0.0375882
rPAD/6182 PAD:5459 PAD:11167 1.5
rPAD/6183 PAD:5458 PAD:5461 0.0375882
rPAD/6184 PAD:5458 PAD:5459 1.5
rPAD/6185 PAD:5456 PAD:5459 0.0751765
rPAD/6186 PAD:5456 PAD:11164 1.5
rPAD/6187 PAD:5455 PAD:5458 0.0751765
rPAD/6188 PAD:5455 PAD:5456 1.5
rPAD/6189 PAD:5453 PAD:5456 0.0375882
rPAD/6190 PAD:5453 PAD:11161 1.5
rPAD/6191 PAD:5452 PAD:5455 0.0375882
rPAD/6192 PAD:5452 PAD:5453 1.5
rPAD/6193 PAD:5450 PAD:5453 0.0751765
rPAD/6194 PAD:5450 PAD:11158 1.5
rPAD/6195 PAD:5449 PAD:5452 0.0751765
rPAD/6196 PAD:5449 PAD:5450 1.5
rPAD/6197 PAD:5447 PAD:11151 0.0751765
rPAD/6198 PAD:5447 PAD:5450 0.0375882
rPAD/6199 PAD:5447 PAD:11155 1.5
rPAD/6200 PAD:5446 PAD:5449 0.0375882
rPAD/6201 PAD:5446 PAD:5447 1.5
rPAD/6202 PAD:5443 PAD:5446 0.0751765
rPAD/6203 PAD:5443 PAD:11151 1.5
rPAD/6204 PAD:5441 PAD:11145 0.0751765
rPAD/6205 PAD:5441 PAD:11151 0.0375882
rPAD/6206 PAD:5441 PAD:11149 1.5
rPAD/6207 PAD:5440 PAD:5443 0.0375882
rPAD/6208 PAD:5440 PAD:5441 1.5
rPAD/6209 PAD:5437 PAD:5440 0.0751765
rPAD/6210 PAD:5437 PAD:11145 1.5
rPAD/6211 PAD:5434 PAD:5437 0.0375882
rPAD/6212 PAD:5434 PAD:11142 1.5
rPAD/6213 PAD:5431 PAD:5434 0.0751765
rPAD/6214 PAD:5431 PAD:11139 1.5
rPAD/6215 PAD:5429 PAD:11133 0.0751765
rPAD/6216 PAD:5429 PAD:11139 0.0375882
rPAD/6217 PAD:5429 PAD:11137 1.5
rPAD/6218 PAD:5428 PAD:5431 0.0375882
rPAD/6219 PAD:5428 PAD:5429 1.5
rPAD/6220 PAD:5425 PAD:5428 0.0751765
rPAD/6221 PAD:5425 PAD:11133 1.5
rPAD/6222 PAD:5422 PAD:5425 0.0375882
rPAD/6223 PAD:5422 PAD:11130 1.5
rPAD/6224 PAD:5420 PAD:11130 0.0751765
rPAD/6225 PAD:5420 PAD:11128 1.5
rPAD/6226 PAD:5419 PAD:5422 0.0751765
rPAD/6227 PAD:5419 PAD:5420 1.5
rPAD/6228 PAD:5417 PAD:5420 0.0375882
rPAD/6229 PAD:5417 PAD:11125 1.5
rPAD/6230 PAD:5416 PAD:5419 0.0375882
rPAD/6231 PAD:5416 PAD:5417 1.5
rPAD/6232 PAD:5414 PAD:5417 0.0751765
rPAD/6233 PAD:5414 PAD:11122 1.5
rPAD/6234 PAD:5413 PAD:5416 0.0751765
rPAD/6235 PAD:5413 PAD:5414 1.5
rPAD/6236 PAD:5411 PAD:5414 0.0375882
rPAD/6237 PAD:5411 PAD:11119 1.5
rPAD/6238 PAD:5410 PAD:5413 0.0375882
rPAD/6239 PAD:5410 PAD:5411 1.5
rPAD/6240 PAD:5408 PAD:5411 0.0751765
rPAD/6241 PAD:5408 PAD:11116 1.5
rPAD/6242 PAD:5407 PAD:5410 0.0751765
rPAD/6243 PAD:5407 PAD:5408 1.5
rPAD/6244 PAD:5405 PAD:11109 0.0751765
rPAD/6245 PAD:5405 PAD:5408 0.0375882
rPAD/6246 PAD:5405 PAD:11113 1.5
rPAD/6247 PAD:5404 PAD:5407 0.0375882
rPAD/6248 PAD:5404 PAD:5405 1.5
rPAD/6249 PAD:5401 PAD:5404 0.0751765
rPAD/6250 PAD:5401 PAD:11109 1.5
rPAD/6251 PAD:5399 PAD:11109 0.0375882
rPAD/6252 PAD:5399 PAD:11107 1.5
rPAD/6253 PAD:5398 PAD:5401 0.0375882
rPAD/6254 PAD:5398 PAD:5399 1.5
rPAD/6255 PAD:5396 PAD:5399 0.0751765
rPAD/6256 PAD:5396 PAD:11104 1.5
rPAD/6257 PAD:5395 PAD:5398 0.0751765
rPAD/6258 PAD:5395 PAD:5396 1.5
rPAD/6259 PAD:5393 PAD:11097 0.0751765
rPAD/6260 PAD:5393 PAD:5396 0.0375882
rPAD/6261 PAD:5393 PAD:11101 1.5
rPAD/6262 PAD:5392 PAD:5395 0.0375882
rPAD/6263 PAD:5392 PAD:5393 1.5
rPAD/6264 PAD:5389 PAD:5392 0.0751765
rPAD/6265 PAD:5389 PAD:11097 1.5
rPAD/6266 PAD:5386 PAD:5389 0.0375882
rPAD/6267 PAD:5386 PAD:11094 1.5
rPAD/6268 PAD:5383 PAD:5386 0.0751765
rPAD/6269 PAD:5383 PAD:11091 1.5
rPAD/6270 PAD:5380 PAD:5383 0.0375882
rPAD/6271 PAD:5380 PAD:11088 1.5
rPAD/6272 PAD:5377 PAD:5380 0.0751765
rPAD/6273 PAD:5377 PAD:11085 1.5
rPAD/6274 PAD:5375 PAD:11085 0.0375882
rPAD/6275 PAD:5375 PAD:11083 1.5
rPAD/6276 PAD:5374 PAD:5377 0.0375882
rPAD/6277 PAD:5374 PAD:5375 1.5
rPAD/6278 PAD:5372 PAD:11076 0.0375882
rPAD/6279 PAD:5372 PAD:5375 0.0751765
rPAD/6280 PAD:5372 PAD:11080 1.5
rPAD/6281 PAD:5371 PAD:5374 0.0751765
rPAD/6282 PAD:5371 PAD:5372 1.5
rPAD/6283 PAD:5368 PAD:5371 0.0375882
rPAD/6284 PAD:5368 PAD:11076 1.5
rPAD/6285 PAD:5366 PAD:11076 0.0751765
rPAD/6286 PAD:5366 PAD:11074 1.5
rPAD/6287 PAD:5365 PAD:5368 0.0751765
rPAD/6288 PAD:5365 PAD:5366 1.5
rPAD/6289 PAD:5363 PAD:5366 0.0375882
rPAD/6290 PAD:5363 PAD:11071 1.5
rPAD/6291 PAD:5362 PAD:5365 0.0375882
rPAD/6292 PAD:5362 PAD:5363 1.5
rPAD/6293 PAD:5360 PAD:5363 0.0751765
rPAD/6294 PAD:5360 PAD:11068 1.5
rPAD/6295 PAD:5359 PAD:5362 0.0751765
rPAD/6296 PAD:5359 PAD:5360 1.5
rPAD/6297 PAD:5357 PAD:5360 0.0375882
rPAD/6298 PAD:5357 PAD:11065 1.5
rPAD/6299 PAD:5356 PAD:5359 0.0375882
rPAD/6300 PAD:5356 PAD:5357 1.5
rPAD/6301 PAD:5354 PAD:5357 0.0751765
rPAD/6302 PAD:5354 PAD:11062 1.5
rPAD/6303 PAD:5353 PAD:5356 0.0751765
rPAD/6304 PAD:5353 PAD:5354 1.5
rPAD/6305 PAD:5351 PAD:11055 0.0751765
rPAD/6306 PAD:5351 PAD:5354 0.0375882
rPAD/6307 PAD:5351 PAD:11059 1.5
rPAD/6308 PAD:5350 PAD:5353 0.0375882
rPAD/6309 PAD:5350 PAD:5351 1.5
rPAD/6310 PAD:5347 PAD:5350 0.0751765
rPAD/6311 PAD:5347 PAD:11055 1.5
rPAD/6312 PAD:5345 PAD:11055 0.0375882
rPAD/6313 PAD:5345 PAD:11053 1.5
rPAD/6314 PAD:5344 PAD:5347 0.0375882
rPAD/6315 PAD:5344 PAD:5345 1.5
rPAD/6316 PAD:5342 PAD:5345 0.0751765
rPAD/6317 PAD:5342 PAD:11050 1.5
rPAD/6318 PAD:5341 PAD:5344 0.0751765
rPAD/6319 PAD:5341 PAD:5342 1.5
rPAD/6320 PAD:5339 PAD:5342 0.0375882
rPAD/6321 PAD:5339 PAD:11047 1.5
rPAD/6322 PAD:5338 PAD:5341 0.0375882
rPAD/6323 PAD:5338 PAD:5339 1.5
rPAD/6324 PAD:5336 PAD:5339 0.0751765
rPAD/6325 PAD:5336 PAD:11044 1.5
rPAD/6326 PAD:5335 PAD:5338 0.0751765
rPAD/6327 PAD:5335 PAD:5336 1.5
rPAD/6328 PAD:5333 PAD:5336 0.0375882
rPAD/6329 PAD:5333 PAD:11041 1.5
rPAD/6330 PAD:5332 PAD:5335 0.0375882
rPAD/6331 PAD:5332 PAD:5333 1.5
rPAD/6332 PAD:5330 PAD:5333 0.0751765
rPAD/6333 PAD:5330 PAD:11038 1.5
rPAD/6334 PAD:5329 PAD:5332 0.0751765
rPAD/6335 PAD:5329 PAD:5330 1.5
rPAD/6336 PAD:5327 PAD:5330 0.0375882
rPAD/6337 PAD:5327 PAD:11035 1.5
rPAD/6338 PAD:5326 PAD:5329 0.0375882
rPAD/6339 PAD:5326 PAD:5327 1.5
rPAD/6340 PAD:5324 PAD:14878 0.0283817
rPAD/6341 PAD:5324 PAD:5327 0.0751765
rPAD/6342 PAD:5324 PAD:11032 1.5
rPAD/6343 PAD:5323 PAD:9157 0.0378785
rPAD/6344 PAD:5323 PAD:5326 0.0751765
rPAD/6345 PAD:5323 PAD:5324 1.5
rPAD/6346 PAD:5319 PAD:10859 0.0100588
rPAD/6347 PAD:5319 PAD:11027 1.5
rPAD/6348 PAD:5318 PAD:9349 0.0670908
rPAD/6349 PAD:5318 PAD:5319 1.5
rPAD/6350 PAD:5316 PAD:5319 0.0751765
rPAD/6351 PAD:5316 PAD:11024 1.5
rPAD/6352 PAD:5315 PAD:5318 0.0751765
rPAD/6353 PAD:5315 PAD:5316 1.5
rPAD/6354 PAD:5313 PAD:11017 0.0751765
rPAD/6355 PAD:5313 PAD:5316 0.0375882
rPAD/6356 PAD:5313 PAD:11021 1.5
rPAD/6357 PAD:5312 PAD:5315 0.0375882
rPAD/6358 PAD:5312 PAD:5313 1.5
rPAD/6359 PAD:5309 PAD:5312 0.0751765
rPAD/6360 PAD:5309 PAD:11017 1.5
rPAD/6361 PAD:5307 PAD:11017 0.0375882
rPAD/6362 PAD:5307 PAD:11015 1.5
rPAD/6363 PAD:5306 PAD:5309 0.0375882
rPAD/6364 PAD:5306 PAD:5307 1.5
rPAD/6365 PAD:5304 PAD:5307 0.0751765
rPAD/6366 PAD:5304 PAD:11012 1.5
rPAD/6367 PAD:5303 PAD:5306 0.0751765
rPAD/6368 PAD:5303 PAD:5304 1.5
rPAD/6369 PAD:5301 PAD:5304 0.0375882
rPAD/6370 PAD:5301 PAD:11009 1.5
rPAD/6371 PAD:5300 PAD:5303 0.0375882
rPAD/6372 PAD:5300 PAD:5301 1.5
rPAD/6373 PAD:5298 PAD:5301 0.0751765
rPAD/6374 PAD:5298 PAD:11006 1.5
rPAD/6375 PAD:5297 PAD:5300 0.0751765
rPAD/6376 PAD:5297 PAD:5298 1.5
rPAD/6377 PAD:5295 PAD:5298 0.0375882
rPAD/6378 PAD:5295 PAD:11003 1.5
rPAD/6379 PAD:5294 PAD:5297 0.0375882
rPAD/6380 PAD:5294 PAD:5295 1.5
rPAD/6381 PAD:5292 PAD:5295 0.0751765
rPAD/6382 PAD:5292 PAD:11000 1.5
rPAD/6383 PAD:5291 PAD:5294 0.0751765
rPAD/6384 PAD:5291 PAD:5292 1.5
rPAD/6385 PAD:5289 PAD:5292 0.0375882
rPAD/6386 PAD:5289 PAD:10997 1.5
rPAD/6387 PAD:5288 PAD:5291 0.0375882
rPAD/6388 PAD:5288 PAD:5289 1.5
rPAD/6389 PAD:5286 PAD:5289 0.0751765
rPAD/6390 PAD:5286 PAD:10994 1.5
rPAD/6391 PAD:5285 PAD:5288 0.0751765
rPAD/6392 PAD:5285 PAD:5286 1.5
rPAD/6393 PAD:5283 PAD:5286 0.0375882
rPAD/6394 PAD:5283 PAD:10991 1.5
rPAD/6395 PAD:5282 PAD:5285 0.0375882
rPAD/6396 PAD:5282 PAD:5283 1.5
rPAD/6397 PAD:5280 PAD:5283 0.0751765
rPAD/6398 PAD:5280 PAD:10988 1.5
rPAD/6399 PAD:5279 PAD:5282 0.0751765
rPAD/6400 PAD:5279 PAD:5280 1.5
rPAD/6401 PAD:5277 PAD:10981 0.0751765
rPAD/6402 PAD:5277 PAD:5280 0.0375882
rPAD/6403 PAD:5277 PAD:10985 1.5
rPAD/6404 PAD:5276 PAD:5279 0.0375882
rPAD/6405 PAD:5276 PAD:5277 1.5
rPAD/6406 PAD:5273 PAD:5276 0.0751765
rPAD/6407 PAD:5273 PAD:10981 1.5
rPAD/6408 PAD:5271 PAD:10975 0.0751765
rPAD/6409 PAD:5271 PAD:10981 0.0375882
rPAD/6410 PAD:5271 PAD:10979 1.5
rPAD/6411 PAD:5270 PAD:5273 0.0375882
rPAD/6412 PAD:5270 PAD:5271 1.5
rPAD/6413 PAD:5267 PAD:5270 0.0751765
rPAD/6414 PAD:5267 PAD:10975 1.5
rPAD/6415 PAD:5264 PAD:5267 0.0375882
rPAD/6416 PAD:5264 PAD:10972 1.5
rPAD/6417 PAD:5261 PAD:5264 0.0751765
rPAD/6418 PAD:5261 PAD:10969 1.5
rPAD/6419 PAD:5259 PAD:10963 0.0751765
rPAD/6420 PAD:5259 PAD:10969 0.0375882
rPAD/6421 PAD:5259 PAD:10967 1.5
rPAD/6422 PAD:5258 PAD:5261 0.0375882
rPAD/6423 PAD:5258 PAD:5259 1.5
rPAD/6424 PAD:5255 PAD:5258 0.0751765
rPAD/6425 PAD:5255 PAD:10963 1.5
rPAD/6426 PAD:5252 PAD:5255 0.0375882
rPAD/6427 PAD:5252 PAD:10960 1.5
rPAD/6428 PAD:5250 PAD:10960 0.0751765
rPAD/6429 PAD:5250 PAD:10958 1.5
rPAD/6430 PAD:5249 PAD:5252 0.0751765
rPAD/6431 PAD:5249 PAD:5250 1.5
rPAD/6432 PAD:5247 PAD:5250 0.0375882
rPAD/6433 PAD:5247 PAD:10955 1.5
rPAD/6434 PAD:5246 PAD:5249 0.0375882
rPAD/6435 PAD:5246 PAD:5247 1.5
rPAD/6436 PAD:5244 PAD:5247 0.0751765
rPAD/6437 PAD:5244 PAD:10952 1.5
rPAD/6438 PAD:5243 PAD:5246 0.0751765
rPAD/6439 PAD:5243 PAD:5244 1.5
rPAD/6440 PAD:5241 PAD:5244 0.0375882
rPAD/6441 PAD:5241 PAD:10949 1.5
rPAD/6442 PAD:5240 PAD:5243 0.0375882
rPAD/6443 PAD:5240 PAD:5241 1.5
rPAD/6444 PAD:5238 PAD:5241 0.0751765
rPAD/6445 PAD:5238 PAD:10946 1.5
rPAD/6446 PAD:5237 PAD:5240 0.0751765
rPAD/6447 PAD:5237 PAD:5238 1.5
rPAD/6448 PAD:5235 PAD:10939 0.0751765
rPAD/6449 PAD:5235 PAD:5238 0.0375882
rPAD/6450 PAD:5235 PAD:10943 1.5
rPAD/6451 PAD:5234 PAD:5237 0.0375882
rPAD/6452 PAD:5234 PAD:5235 1.5
rPAD/6453 PAD:5231 PAD:5234 0.0751765
rPAD/6454 PAD:5231 PAD:10939 1.5
rPAD/6455 PAD:5229 PAD:10939 0.0375882
rPAD/6456 PAD:5229 PAD:10937 1.5
rPAD/6457 PAD:5228 PAD:5231 0.0375882
rPAD/6458 PAD:5228 PAD:5229 1.5
rPAD/6459 PAD:5226 PAD:5229 0.0751765
rPAD/6460 PAD:5226 PAD:10934 1.5
rPAD/6461 PAD:5225 PAD:5228 0.0751765
rPAD/6462 PAD:5225 PAD:5226 1.5
rPAD/6463 PAD:5223 PAD:10927 0.0751765
rPAD/6464 PAD:5223 PAD:5226 0.0375882
rPAD/6465 PAD:5223 PAD:10931 1.5
rPAD/6466 PAD:5222 PAD:5225 0.0375882
rPAD/6467 PAD:5222 PAD:5223 1.5
rPAD/6468 PAD:5219 PAD:5222 0.0751765
rPAD/6469 PAD:5219 PAD:10927 1.5
rPAD/6470 PAD:5216 PAD:5219 0.0375882
rPAD/6471 PAD:5216 PAD:10924 1.5
rPAD/6472 PAD:5213 PAD:5216 0.0751765
rPAD/6473 PAD:5213 PAD:10921 1.5
rPAD/6474 PAD:5210 PAD:5213 0.0375882
rPAD/6475 PAD:5210 PAD:10918 1.5
rPAD/6476 PAD:5207 PAD:5210 0.0751765
rPAD/6477 PAD:5207 PAD:10915 1.5
rPAD/6478 PAD:5205 PAD:10915 0.0375882
rPAD/6479 PAD:5205 PAD:10913 1.5
rPAD/6480 PAD:5204 PAD:5207 0.0375882
rPAD/6481 PAD:5204 PAD:5205 1.5
rPAD/6482 PAD:5202 PAD:10906 0.0375882
rPAD/6483 PAD:5202 PAD:5205 0.0751765
rPAD/6484 PAD:5202 PAD:10910 1.5
rPAD/6485 PAD:5201 PAD:5204 0.0751765
rPAD/6486 PAD:5201 PAD:5202 1.5
rPAD/6487 PAD:5198 PAD:5201 0.0375882
rPAD/6488 PAD:5198 PAD:10906 1.5
rPAD/6489 PAD:5196 PAD:10906 0.0751765
rPAD/6490 PAD:5196 PAD:10904 1.5
rPAD/6491 PAD:5195 PAD:5198 0.0751765
rPAD/6492 PAD:5195 PAD:5196 1.5
rPAD/6493 PAD:5193 PAD:5196 0.0375882
rPAD/6494 PAD:5193 PAD:10901 1.5
rPAD/6495 PAD:5192 PAD:5195 0.0375882
rPAD/6496 PAD:5192 PAD:5193 1.5
rPAD/6497 PAD:5190 PAD:5193 0.0751765
rPAD/6498 PAD:5190 PAD:10898 1.5
rPAD/6499 PAD:5189 PAD:5192 0.0751765
rPAD/6500 PAD:5189 PAD:5190 1.5
rPAD/6501 PAD:5187 PAD:5190 0.0375882
rPAD/6502 PAD:5187 PAD:10895 1.5
rPAD/6503 PAD:5186 PAD:5189 0.0375882
rPAD/6504 PAD:5186 PAD:5187 1.5
rPAD/6505 PAD:5184 PAD:5187 0.0751765
rPAD/6506 PAD:5184 PAD:10892 1.5
rPAD/6507 PAD:5183 PAD:5186 0.0751765
rPAD/6508 PAD:5183 PAD:5184 1.5
rPAD/6509 PAD:5181 PAD:10885 0.0751765
rPAD/6510 PAD:5181 PAD:5184 0.0375882
rPAD/6511 PAD:5181 PAD:10889 1.5
rPAD/6512 PAD:5180 PAD:5183 0.0375882
rPAD/6513 PAD:5180 PAD:5181 1.5
rPAD/6514 PAD:5177 PAD:5180 0.0751765
rPAD/6515 PAD:5177 PAD:10885 1.5
rPAD/6516 PAD:5175 PAD:10885 0.0375882
rPAD/6517 PAD:5175 PAD:10883 1.5
rPAD/6518 PAD:5174 PAD:5177 0.0375882
rPAD/6519 PAD:5174 PAD:5175 1.5
rPAD/6520 PAD:5172 PAD:5175 0.0751765
rPAD/6521 PAD:5172 PAD:10880 1.5
rPAD/6522 PAD:5171 PAD:5174 0.0751765
rPAD/6523 PAD:5171 PAD:5172 1.5
rPAD/6524 PAD:5169 PAD:5172 0.0375882
rPAD/6525 PAD:5169 PAD:10877 1.5
rPAD/6526 PAD:5168 PAD:5171 0.0375882
rPAD/6527 PAD:5168 PAD:5169 1.5
rPAD/6528 PAD:5166 PAD:5169 0.0751765
rPAD/6529 PAD:5166 PAD:10874 1.5
rPAD/6530 PAD:5165 PAD:5168 0.0751765
rPAD/6531 PAD:5165 PAD:5166 1.5
rPAD/6532 PAD:5163 PAD:5166 0.0375882
rPAD/6533 PAD:5163 PAD:10871 1.5
rPAD/6534 PAD:5162 PAD:5165 0.0375882
rPAD/6535 PAD:5162 PAD:5163 1.5
rPAD/6536 PAD:5160 PAD:5163 0.0751765
rPAD/6537 PAD:5160 PAD:10868 1.5
rPAD/6538 PAD:5159 PAD:5162 0.0751765
rPAD/6539 PAD:5159 PAD:5160 1.5
rPAD/6540 PAD:5157 PAD:5160 0.0375882
rPAD/6541 PAD:5157 PAD:10865 1.5
rPAD/6542 PAD:5156 PAD:5159 0.0375882
rPAD/6543 PAD:5156 PAD:5157 1.5
rPAD/6544 PAD:5154 PAD:14873 0.0283817
rPAD/6545 PAD:5154 PAD:5157 0.0751765
rPAD/6546 PAD:5154 PAD:10862 1.5
rPAD/6547 PAD:5153 PAD:9150 0.0378785
rPAD/6548 PAD:5153 PAD:5156 0.0751765
rPAD/6549 PAD:5153 PAD:5154 1.5
rPAD/6550 PAD:5149 PAD:10689 0.0100588
rPAD/6551 PAD:5149 PAD:10857 1.5
rPAD/6552 PAD:5148 PAD:9344 0.0670908
rPAD/6553 PAD:5148 PAD:5149 1.5
rPAD/6554 PAD:5146 PAD:5149 0.0751765
rPAD/6555 PAD:5146 PAD:10854 1.5
rPAD/6556 PAD:5145 PAD:5148 0.0751765
rPAD/6557 PAD:5145 PAD:5146 1.5
rPAD/6558 PAD:5143 PAD:10847 0.0751765
rPAD/6559 PAD:5143 PAD:5146 0.0375882
rPAD/6560 PAD:5143 PAD:10851 1.5
rPAD/6561 PAD:5142 PAD:5145 0.0375882
rPAD/6562 PAD:5142 PAD:5143 1.5
rPAD/6563 PAD:5139 PAD:5142 0.0751765
rPAD/6564 PAD:5139 PAD:10847 1.5
rPAD/6565 PAD:5137 PAD:10847 0.0375882
rPAD/6566 PAD:5137 PAD:10845 1.5
rPAD/6567 PAD:5136 PAD:5139 0.0375882
rPAD/6568 PAD:5136 PAD:5137 1.5
rPAD/6569 PAD:5134 PAD:5137 0.0751765
rPAD/6570 PAD:5134 PAD:10842 1.5
rPAD/6571 PAD:5133 PAD:5136 0.0751765
rPAD/6572 PAD:5133 PAD:5134 1.5
rPAD/6573 PAD:5131 PAD:5134 0.0375882
rPAD/6574 PAD:5131 PAD:10839 1.5
rPAD/6575 PAD:5130 PAD:5133 0.0375882
rPAD/6576 PAD:5130 PAD:5131 1.5
rPAD/6577 PAD:5128 PAD:5131 0.0751765
rPAD/6578 PAD:5128 PAD:10836 1.5
rPAD/6579 PAD:5127 PAD:5130 0.0751765
rPAD/6580 PAD:5127 PAD:5128 1.5
rPAD/6581 PAD:5125 PAD:5128 0.0375882
rPAD/6582 PAD:5125 PAD:10833 1.5
rPAD/6583 PAD:5124 PAD:5127 0.0375882
rPAD/6584 PAD:5124 PAD:5125 1.5
rPAD/6585 PAD:5122 PAD:5125 0.0751765
rPAD/6586 PAD:5122 PAD:10830 1.5
rPAD/6587 PAD:5121 PAD:5124 0.0751765
rPAD/6588 PAD:5121 PAD:5122 1.5
rPAD/6589 PAD:5119 PAD:5122 0.0375882
rPAD/6590 PAD:5119 PAD:10827 1.5
rPAD/6591 PAD:5118 PAD:5121 0.0375882
rPAD/6592 PAD:5118 PAD:5119 1.5
rPAD/6593 PAD:5116 PAD:5119 0.0751765
rPAD/6594 PAD:5116 PAD:10824 1.5
rPAD/6595 PAD:5115 PAD:5118 0.0751765
rPAD/6596 PAD:5115 PAD:5116 1.5
rPAD/6597 PAD:5113 PAD:5116 0.0375882
rPAD/6598 PAD:5113 PAD:10821 1.5
rPAD/6599 PAD:5112 PAD:5115 0.0375882
rPAD/6600 PAD:5112 PAD:5113 1.5
rPAD/6601 PAD:5110 PAD:5113 0.0751765
rPAD/6602 PAD:5110 PAD:10818 1.5
rPAD/6603 PAD:5109 PAD:5112 0.0751765
rPAD/6604 PAD:5109 PAD:5110 1.5
rPAD/6605 PAD:5107 PAD:10811 0.0751765
rPAD/6606 PAD:5107 PAD:5110 0.0375882
rPAD/6607 PAD:5107 PAD:10815 1.5
rPAD/6608 PAD:5106 PAD:5109 0.0375882
rPAD/6609 PAD:5106 PAD:5107 1.5
rPAD/6610 PAD:5103 PAD:5106 0.0751765
rPAD/6611 PAD:5103 PAD:10811 1.5
rPAD/6612 PAD:5101 PAD:10805 0.0751765
rPAD/6613 PAD:5101 PAD:10811 0.0375882
rPAD/6614 PAD:5101 PAD:10809 1.5
rPAD/6615 PAD:5100 PAD:5103 0.0375882
rPAD/6616 PAD:5100 PAD:5101 1.5
rPAD/6617 PAD:5097 PAD:5100 0.0751765
rPAD/6618 PAD:5097 PAD:10805 1.5
rPAD/6619 PAD:5094 PAD:5097 0.0375882
rPAD/6620 PAD:5094 PAD:10802 1.5
rPAD/6621 PAD:5091 PAD:5094 0.0751765
rPAD/6622 PAD:5091 PAD:10799 1.5
rPAD/6623 PAD:5089 PAD:10793 0.0751765
rPAD/6624 PAD:5089 PAD:10799 0.0375882
rPAD/6625 PAD:5089 PAD:10797 1.5
rPAD/6626 PAD:5088 PAD:5091 0.0375882
rPAD/6627 PAD:5088 PAD:5089 1.5
rPAD/6628 PAD:5085 PAD:5088 0.0751765
rPAD/6629 PAD:5085 PAD:10793 1.5
rPAD/6630 PAD:5082 PAD:5085 0.0375882
rPAD/6631 PAD:5082 PAD:10790 1.5
rPAD/6632 PAD:5080 PAD:10790 0.0751765
rPAD/6633 PAD:5080 PAD:10788 1.5
rPAD/6634 PAD:5079 PAD:5082 0.0751765
rPAD/6635 PAD:5079 PAD:5080 1.5
rPAD/6636 PAD:5077 PAD:5080 0.0375882
rPAD/6637 PAD:5077 PAD:10785 1.5
rPAD/6638 PAD:5076 PAD:5079 0.0375882
rPAD/6639 PAD:5076 PAD:5077 1.5
rPAD/6640 PAD:5074 PAD:5077 0.0751765
rPAD/6641 PAD:5074 PAD:10782 1.5
rPAD/6642 PAD:5073 PAD:5076 0.0751765
rPAD/6643 PAD:5073 PAD:5074 1.5
rPAD/6644 PAD:5071 PAD:5074 0.0375882
rPAD/6645 PAD:5071 PAD:10779 1.5
rPAD/6646 PAD:5070 PAD:5073 0.0375882
rPAD/6647 PAD:5070 PAD:5071 1.5
rPAD/6648 PAD:5068 PAD:5071 0.0751765
rPAD/6649 PAD:5068 PAD:10776 1.5
rPAD/6650 PAD:5067 PAD:5070 0.0751765
rPAD/6651 PAD:5067 PAD:5068 1.5
rPAD/6652 PAD:5065 PAD:10769 0.0751765
rPAD/6653 PAD:5065 PAD:5068 0.0375882
rPAD/6654 PAD:5065 PAD:10773 1.5
rPAD/6655 PAD:5064 PAD:5067 0.0375882
rPAD/6656 PAD:5064 PAD:5065 1.5
rPAD/6657 PAD:5061 PAD:5064 0.0751765
rPAD/6658 PAD:5061 PAD:10769 1.5
rPAD/6659 PAD:5059 PAD:10769 0.0375882
rPAD/6660 PAD:5059 PAD:10767 1.5
rPAD/6661 PAD:5058 PAD:5061 0.0375882
rPAD/6662 PAD:5058 PAD:5059 1.5
rPAD/6663 PAD:5056 PAD:5059 0.0751765
rPAD/6664 PAD:5056 PAD:10764 1.5
rPAD/6665 PAD:5055 PAD:5058 0.0751765
rPAD/6666 PAD:5055 PAD:5056 1.5
rPAD/6667 PAD:5053 PAD:10757 0.0751765
rPAD/6668 PAD:5053 PAD:5056 0.0375882
rPAD/6669 PAD:5053 PAD:10761 1.5
rPAD/6670 PAD:5052 PAD:5055 0.0375882
rPAD/6671 PAD:5052 PAD:5053 1.5
rPAD/6672 PAD:5049 PAD:5052 0.0751765
rPAD/6673 PAD:5049 PAD:10757 1.5
rPAD/6674 PAD:5046 PAD:5049 0.0375882
rPAD/6675 PAD:5046 PAD:10754 1.5
rPAD/6676 PAD:5043 PAD:5046 0.0751765
rPAD/6677 PAD:5043 PAD:10751 1.5
rPAD/6678 PAD:5040 PAD:5043 0.0375882
rPAD/6679 PAD:5040 PAD:10748 1.5
rPAD/6680 PAD:5037 PAD:5040 0.0751765
rPAD/6681 PAD:5037 PAD:10745 1.5
rPAD/6682 PAD:5035 PAD:10745 0.0375882
rPAD/6683 PAD:5035 PAD:10743 1.5
rPAD/6684 PAD:5034 PAD:5037 0.0375882
rPAD/6685 PAD:5034 PAD:5035 1.5
rPAD/6686 PAD:5032 PAD:10736 0.0375882
rPAD/6687 PAD:5032 PAD:5035 0.0751765
rPAD/6688 PAD:5032 PAD:10740 1.5
rPAD/6689 PAD:5031 PAD:5034 0.0751765
rPAD/6690 PAD:5031 PAD:5032 1.5
rPAD/6691 PAD:5028 PAD:5031 0.0375882
rPAD/6692 PAD:5028 PAD:10736 1.5
rPAD/6693 PAD:5026 PAD:10736 0.0751765
rPAD/6694 PAD:5026 PAD:10734 1.5
rPAD/6695 PAD:5025 PAD:5028 0.0751765
rPAD/6696 PAD:5025 PAD:5026 1.5
rPAD/6697 PAD:5023 PAD:5026 0.0375882
rPAD/6698 PAD:5023 PAD:10731 1.5
rPAD/6699 PAD:5022 PAD:5025 0.0375882
rPAD/6700 PAD:5022 PAD:5023 1.5
rPAD/6701 PAD:5020 PAD:5023 0.0751765
rPAD/6702 PAD:5020 PAD:10728 1.5
rPAD/6703 PAD:5019 PAD:5022 0.0751765
rPAD/6704 PAD:5019 PAD:5020 1.5
rPAD/6705 PAD:5017 PAD:5020 0.0375882
rPAD/6706 PAD:5017 PAD:10725 1.5
rPAD/6707 PAD:5016 PAD:5019 0.0375882
rPAD/6708 PAD:5016 PAD:5017 1.5
rPAD/6709 PAD:5014 PAD:5017 0.0751765
rPAD/6710 PAD:5014 PAD:10722 1.5
rPAD/6711 PAD:5013 PAD:5016 0.0751765
rPAD/6712 PAD:5013 PAD:5014 1.5
rPAD/6713 PAD:5011 PAD:10715 0.0751765
rPAD/6714 PAD:5011 PAD:5014 0.0375882
rPAD/6715 PAD:5011 PAD:10719 1.5
rPAD/6716 PAD:5010 PAD:5013 0.0375882
rPAD/6717 PAD:5010 PAD:5011 1.5
rPAD/6718 PAD:5007 PAD:5010 0.0751765
rPAD/6719 PAD:5007 PAD:10715 1.5
rPAD/6720 PAD:5005 PAD:10715 0.0375882
rPAD/6721 PAD:5005 PAD:10713 1.5
rPAD/6722 PAD:5004 PAD:5007 0.0375882
rPAD/6723 PAD:5004 PAD:5005 1.5
rPAD/6724 PAD:5002 PAD:5005 0.0751765
rPAD/6725 PAD:5002 PAD:10710 1.5
rPAD/6726 PAD:5001 PAD:5004 0.0751765
rPAD/6727 PAD:5001 PAD:5002 1.5
rPAD/6728 PAD:4999 PAD:5002 0.0375882
rPAD/6729 PAD:4999 PAD:10707 1.5
rPAD/6730 PAD:4998 PAD:5001 0.0375882
rPAD/6731 PAD:4998 PAD:4999 1.5
rPAD/6732 PAD:4996 PAD:4999 0.0751765
rPAD/6733 PAD:4996 PAD:10704 1.5
rPAD/6734 PAD:4995 PAD:4998 0.0751765
rPAD/6735 PAD:4995 PAD:4996 1.5
rPAD/6736 PAD:4993 PAD:4996 0.0375882
rPAD/6737 PAD:4993 PAD:10701 1.5
rPAD/6738 PAD:4992 PAD:4995 0.0375882
rPAD/6739 PAD:4992 PAD:4993 1.5
rPAD/6740 PAD:4990 PAD:4993 0.0751765
rPAD/6741 PAD:4990 PAD:10698 1.5
rPAD/6742 PAD:4989 PAD:4992 0.0751765
rPAD/6743 PAD:4989 PAD:4990 1.5
rPAD/6744 PAD:4987 PAD:4990 0.0375882
rPAD/6745 PAD:4987 PAD:10695 1.5
rPAD/6746 PAD:4986 PAD:4989 0.0375882
rPAD/6747 PAD:4986 PAD:4987 1.5
rPAD/6748 PAD:4984 PAD:14867 0.0283817
rPAD/6749 PAD:4984 PAD:4987 0.0751765
rPAD/6750 PAD:4984 PAD:10692 1.5
rPAD/6751 PAD:4983 PAD:9143 0.0378785
rPAD/6752 PAD:4983 PAD:4986 0.0751765
rPAD/6753 PAD:4983 PAD:4984 1.5
rPAD/6754 PAD:4979 PAD:10519 0.0100588
rPAD/6755 PAD:4979 PAD:10687 1.5
rPAD/6756 PAD:4978 PAD:9340 0.0670908
rPAD/6757 PAD:4978 PAD:4979 1.5
rPAD/6758 PAD:4976 PAD:4979 0.0751765
rPAD/6759 PAD:4976 PAD:10684 1.5
rPAD/6760 PAD:4975 PAD:4978 0.0751765
rPAD/6761 PAD:4975 PAD:4976 1.5
rPAD/6762 PAD:4973 PAD:10677 0.0751765
rPAD/6763 PAD:4973 PAD:4976 0.0375882
rPAD/6764 PAD:4973 PAD:10681 1.5
rPAD/6765 PAD:4972 PAD:4975 0.0375882
rPAD/6766 PAD:4972 PAD:4973 1.5
rPAD/6767 PAD:4969 PAD:4972 0.0751765
rPAD/6768 PAD:4969 PAD:10677 1.5
rPAD/6769 PAD:4967 PAD:10677 0.0375882
rPAD/6770 PAD:4967 PAD:10675 1.5
rPAD/6771 PAD:4966 PAD:4969 0.0375882
rPAD/6772 PAD:4966 PAD:4967 1.5
rPAD/6773 PAD:4964 PAD:4967 0.0751765
rPAD/6774 PAD:4964 PAD:10672 1.5
rPAD/6775 PAD:4963 PAD:4966 0.0751765
rPAD/6776 PAD:4963 PAD:4964 1.5
rPAD/6777 PAD:4961 PAD:4964 0.0375882
rPAD/6778 PAD:4961 PAD:10669 1.5
rPAD/6779 PAD:4960 PAD:4963 0.0375882
rPAD/6780 PAD:4960 PAD:4961 1.5
rPAD/6781 PAD:4958 PAD:4961 0.0751765
rPAD/6782 PAD:4958 PAD:10666 1.5
rPAD/6783 PAD:4957 PAD:4960 0.0751765
rPAD/6784 PAD:4957 PAD:4958 1.5
rPAD/6785 PAD:4955 PAD:4958 0.0375882
rPAD/6786 PAD:4955 PAD:10663 1.5
rPAD/6787 PAD:4954 PAD:4957 0.0375882
rPAD/6788 PAD:4954 PAD:4955 1.5
rPAD/6789 PAD:4952 PAD:4955 0.0751765
rPAD/6790 PAD:4952 PAD:10660 1.5
rPAD/6791 PAD:4951 PAD:4954 0.0751765
rPAD/6792 PAD:4951 PAD:4952 1.5
rPAD/6793 PAD:4949 PAD:4952 0.0375882
rPAD/6794 PAD:4949 PAD:10657 1.5
rPAD/6795 PAD:4948 PAD:4951 0.0375882
rPAD/6796 PAD:4948 PAD:4949 1.5
rPAD/6797 PAD:4946 PAD:4949 0.0751765
rPAD/6798 PAD:4946 PAD:10654 1.5
rPAD/6799 PAD:4945 PAD:4948 0.0751765
rPAD/6800 PAD:4945 PAD:4946 1.5
rPAD/6801 PAD:4943 PAD:4946 0.0375882
rPAD/6802 PAD:4943 PAD:10651 1.5
rPAD/6803 PAD:4942 PAD:4945 0.0375882
rPAD/6804 PAD:4942 PAD:4943 1.5
rPAD/6805 PAD:4940 PAD:4943 0.0751765
rPAD/6806 PAD:4940 PAD:10648 1.5
rPAD/6807 PAD:4939 PAD:4942 0.0751765
rPAD/6808 PAD:4939 PAD:4940 1.5
rPAD/6809 PAD:4937 PAD:10641 0.0751765
rPAD/6810 PAD:4937 PAD:4940 0.0375882
rPAD/6811 PAD:4937 PAD:10645 1.5
rPAD/6812 PAD:4936 PAD:4939 0.0375882
rPAD/6813 PAD:4936 PAD:4937 1.5
rPAD/6814 PAD:4933 PAD:4936 0.0751765
rPAD/6815 PAD:4933 PAD:10641 1.5
rPAD/6816 PAD:4931 PAD:10635 0.0751765
rPAD/6817 PAD:4931 PAD:10641 0.0375882
rPAD/6818 PAD:4931 PAD:10639 1.5
rPAD/6819 PAD:4930 PAD:4933 0.0375882
rPAD/6820 PAD:4930 PAD:4931 1.5
rPAD/6821 PAD:4927 PAD:4930 0.0751765
rPAD/6822 PAD:4927 PAD:10635 1.5
rPAD/6823 PAD:4924 PAD:4927 0.0375882
rPAD/6824 PAD:4924 PAD:10632 1.5
rPAD/6825 PAD:4921 PAD:4924 0.0751765
rPAD/6826 PAD:4921 PAD:10629 1.5
rPAD/6827 PAD:4919 PAD:10623 0.0751765
rPAD/6828 PAD:4919 PAD:10629 0.0375882
rPAD/6829 PAD:4919 PAD:10627 1.5
rPAD/6830 PAD:4918 PAD:4921 0.0375882
rPAD/6831 PAD:4918 PAD:4919 1.5
rPAD/6832 PAD:4915 PAD:4918 0.0751765
rPAD/6833 PAD:4915 PAD:10623 1.5
rPAD/6834 PAD:4912 PAD:4915 0.0375882
rPAD/6835 PAD:4912 PAD:10620 1.5
rPAD/6836 PAD:4910 PAD:10620 0.0751765
rPAD/6837 PAD:4910 PAD:10618 1.5
rPAD/6838 PAD:4909 PAD:4912 0.0751765
rPAD/6839 PAD:4909 PAD:4910 1.5
rPAD/6840 PAD:4907 PAD:4910 0.0375882
rPAD/6841 PAD:4907 PAD:10615 1.5
rPAD/6842 PAD:4906 PAD:4909 0.0375882
rPAD/6843 PAD:4906 PAD:4907 1.5
rPAD/6844 PAD:4904 PAD:4907 0.0751765
rPAD/6845 PAD:4904 PAD:10612 1.5
rPAD/6846 PAD:4903 PAD:4906 0.0751765
rPAD/6847 PAD:4903 PAD:4904 1.5
rPAD/6848 PAD:4901 PAD:4904 0.0375882
rPAD/6849 PAD:4901 PAD:10609 1.5
rPAD/6850 PAD:4900 PAD:4903 0.0375882
rPAD/6851 PAD:4900 PAD:4901 1.5
rPAD/6852 PAD:4898 PAD:4901 0.0751765
rPAD/6853 PAD:4898 PAD:10606 1.5
rPAD/6854 PAD:4897 PAD:4900 0.0751765
rPAD/6855 PAD:4897 PAD:4898 1.5
rPAD/6856 PAD:4895 PAD:10599 0.0751765
rPAD/6857 PAD:4895 PAD:4898 0.0375882
rPAD/6858 PAD:4895 PAD:10603 1.5
rPAD/6859 PAD:4894 PAD:4897 0.0375882
rPAD/6860 PAD:4894 PAD:4895 1.5
rPAD/6861 PAD:4891 PAD:4894 0.0751765
rPAD/6862 PAD:4891 PAD:10599 1.5
rPAD/6863 PAD:4889 PAD:10599 0.0375882
rPAD/6864 PAD:4889 PAD:10597 1.5
rPAD/6865 PAD:4888 PAD:4891 0.0375882
rPAD/6866 PAD:4888 PAD:4889 1.5
rPAD/6867 PAD:4886 PAD:4889 0.0751765
rPAD/6868 PAD:4886 PAD:10594 1.5
rPAD/6869 PAD:4885 PAD:4888 0.0751765
rPAD/6870 PAD:4885 PAD:4886 1.5
rPAD/6871 PAD:4883 PAD:10587 0.0751765
rPAD/6872 PAD:4883 PAD:4886 0.0375882
rPAD/6873 PAD:4883 PAD:10591 1.5
rPAD/6874 PAD:4882 PAD:4885 0.0375882
rPAD/6875 PAD:4882 PAD:4883 1.5
rPAD/6876 PAD:4879 PAD:4882 0.0751765
rPAD/6877 PAD:4879 PAD:10587 1.5
rPAD/6878 PAD:4876 PAD:4879 0.0375882
rPAD/6879 PAD:4876 PAD:10584 1.5
rPAD/6880 PAD:4873 PAD:4876 0.0751765
rPAD/6881 PAD:4873 PAD:10581 1.5
rPAD/6882 PAD:4870 PAD:4873 0.0375882
rPAD/6883 PAD:4870 PAD:10578 1.5
rPAD/6884 PAD:4867 PAD:4870 0.0751765
rPAD/6885 PAD:4867 PAD:10575 1.5
rPAD/6886 PAD:4865 PAD:10575 0.0375882
rPAD/6887 PAD:4865 PAD:10573 1.5
rPAD/6888 PAD:4864 PAD:4867 0.0375882
rPAD/6889 PAD:4864 PAD:4865 1.5
rPAD/6890 PAD:4862 PAD:10566 0.0375882
rPAD/6891 PAD:4862 PAD:4865 0.0751765
rPAD/6892 PAD:4862 PAD:10570 1.5
rPAD/6893 PAD:4861 PAD:4864 0.0751765
rPAD/6894 PAD:4861 PAD:4862 1.5
rPAD/6895 PAD:4858 PAD:4861 0.0375882
rPAD/6896 PAD:4858 PAD:10566 1.5
rPAD/6897 PAD:4856 PAD:10566 0.0751765
rPAD/6898 PAD:4856 PAD:10564 1.5
rPAD/6899 PAD:4855 PAD:4858 0.0751765
rPAD/6900 PAD:4855 PAD:4856 1.5
rPAD/6901 PAD:4853 PAD:4856 0.0375882
rPAD/6902 PAD:4853 PAD:10561 1.5
rPAD/6903 PAD:4852 PAD:4855 0.0375882
rPAD/6904 PAD:4852 PAD:4853 1.5
rPAD/6905 PAD:4850 PAD:4853 0.0751765
rPAD/6906 PAD:4850 PAD:10558 1.5
rPAD/6907 PAD:4849 PAD:4852 0.0751765
rPAD/6908 PAD:4849 PAD:4850 1.5
rPAD/6909 PAD:4847 PAD:4850 0.0375882
rPAD/6910 PAD:4847 PAD:10555 1.5
rPAD/6911 PAD:4846 PAD:4849 0.0375882
rPAD/6912 PAD:4846 PAD:4847 1.5
rPAD/6913 PAD:4844 PAD:4847 0.0751765
rPAD/6914 PAD:4844 PAD:10552 1.5
rPAD/6915 PAD:4843 PAD:4846 0.0751765
rPAD/6916 PAD:4843 PAD:4844 1.5
rPAD/6917 PAD:4841 PAD:10545 0.0751765
rPAD/6918 PAD:4841 PAD:4844 0.0375882
rPAD/6919 PAD:4841 PAD:10549 1.5
rPAD/6920 PAD:4840 PAD:4843 0.0375882
rPAD/6921 PAD:4840 PAD:4841 1.5
rPAD/6922 PAD:4837 PAD:4840 0.0751765
rPAD/6923 PAD:4837 PAD:10545 1.5
rPAD/6924 PAD:4835 PAD:10545 0.0375882
rPAD/6925 PAD:4835 PAD:10543 1.5
rPAD/6926 PAD:4834 PAD:4837 0.0375882
rPAD/6927 PAD:4834 PAD:4835 1.5
rPAD/6928 PAD:4832 PAD:4835 0.0751765
rPAD/6929 PAD:4832 PAD:10540 1.5
rPAD/6930 PAD:4831 PAD:4834 0.0751765
rPAD/6931 PAD:4831 PAD:4832 1.5
rPAD/6932 PAD:4829 PAD:4832 0.0375882
rPAD/6933 PAD:4829 PAD:10537 1.5
rPAD/6934 PAD:4828 PAD:4831 0.0375882
rPAD/6935 PAD:4828 PAD:4829 1.5
rPAD/6936 PAD:4826 PAD:4829 0.0751765
rPAD/6937 PAD:4826 PAD:10534 1.5
rPAD/6938 PAD:4825 PAD:4828 0.0751765
rPAD/6939 PAD:4825 PAD:4826 1.5
rPAD/6940 PAD:4823 PAD:4826 0.0375882
rPAD/6941 PAD:4823 PAD:10531 1.5
rPAD/6942 PAD:4822 PAD:4825 0.0375882
rPAD/6943 PAD:4822 PAD:4823 1.5
rPAD/6944 PAD:4820 PAD:4823 0.0751765
rPAD/6945 PAD:4820 PAD:10528 1.5
rPAD/6946 PAD:4819 PAD:4822 0.0751765
rPAD/6947 PAD:4819 PAD:4820 1.5
rPAD/6948 PAD:4817 PAD:4820 0.0375882
rPAD/6949 PAD:4817 PAD:10525 1.5
rPAD/6950 PAD:4816 PAD:4819 0.0375882
rPAD/6951 PAD:4816 PAD:4817 1.5
rPAD/6952 PAD:4814 PAD:14861 0.0283817
rPAD/6953 PAD:4814 PAD:4817 0.0751765
rPAD/6954 PAD:4814 PAD:10522 1.5
rPAD/6955 PAD:4813 PAD:9136 0.0378785
rPAD/6956 PAD:4813 PAD:4816 0.0751765
rPAD/6957 PAD:4813 PAD:4814 1.5
rPAD/6958 PAD:4809 PAD:10349 0.0100588
rPAD/6959 PAD:4809 PAD:10517 1.5
rPAD/6960 PAD:4808 PAD:9336 0.0670908
rPAD/6961 PAD:4808 PAD:4809 1.5
rPAD/6962 PAD:4806 PAD:4809 0.0751765
rPAD/6963 PAD:4806 PAD:10514 1.5
rPAD/6964 PAD:4805 PAD:4808 0.0751765
rPAD/6965 PAD:4805 PAD:4806 1.5
rPAD/6966 PAD:4803 PAD:10507 0.0751765
rPAD/6967 PAD:4803 PAD:4806 0.0375882
rPAD/6968 PAD:4803 PAD:10511 1.5
rPAD/6969 PAD:4802 PAD:4805 0.0375882
rPAD/6970 PAD:4802 PAD:4803 1.5
rPAD/6971 PAD:4799 PAD:4802 0.0751765
rPAD/6972 PAD:4799 PAD:10507 1.5
rPAD/6973 PAD:4797 PAD:10507 0.0375882
rPAD/6974 PAD:4797 PAD:10505 1.5
rPAD/6975 PAD:4796 PAD:4799 0.0375882
rPAD/6976 PAD:4796 PAD:4797 1.5
rPAD/6977 PAD:4794 PAD:4797 0.0751765
rPAD/6978 PAD:4794 PAD:10502 1.5
rPAD/6979 PAD:4793 PAD:4796 0.0751765
rPAD/6980 PAD:4793 PAD:4794 1.5
rPAD/6981 PAD:4791 PAD:4794 0.0375882
rPAD/6982 PAD:4791 PAD:10499 1.5
rPAD/6983 PAD:4790 PAD:4793 0.0375882
rPAD/6984 PAD:4790 PAD:4791 1.5
rPAD/6985 PAD:4788 PAD:4791 0.0751765
rPAD/6986 PAD:4788 PAD:10496 1.5
rPAD/6987 PAD:4787 PAD:4790 0.0751765
rPAD/6988 PAD:4787 PAD:4788 1.5
rPAD/6989 PAD:4785 PAD:4788 0.0375882
rPAD/6990 PAD:4785 PAD:10493 1.5
rPAD/6991 PAD:4784 PAD:4787 0.0375882
rPAD/6992 PAD:4784 PAD:4785 1.5
rPAD/6993 PAD:4782 PAD:4785 0.0751765
rPAD/6994 PAD:4782 PAD:10490 1.5
rPAD/6995 PAD:4781 PAD:4784 0.0751765
rPAD/6996 PAD:4781 PAD:4782 1.5
rPAD/6997 PAD:4779 PAD:4782 0.0375882
rPAD/6998 PAD:4779 PAD:10487 1.5
rPAD/6999 PAD:4778 PAD:4781 0.0375882
rPAD/7000 PAD:4778 PAD:4779 1.5
rPAD/7001 PAD:4776 PAD:4779 0.0751765
rPAD/7002 PAD:4776 PAD:10484 1.5
rPAD/7003 PAD:4775 PAD:4778 0.0751765
rPAD/7004 PAD:4775 PAD:4776 1.5
rPAD/7005 PAD:4773 PAD:4776 0.0375882
rPAD/7006 PAD:4773 PAD:10481 1.5
rPAD/7007 PAD:4772 PAD:4775 0.0375882
rPAD/7008 PAD:4772 PAD:4773 1.5
rPAD/7009 PAD:4770 PAD:4773 0.0751765
rPAD/7010 PAD:4770 PAD:10478 1.5
rPAD/7011 PAD:4769 PAD:4772 0.0751765
rPAD/7012 PAD:4769 PAD:4770 1.5
rPAD/7013 PAD:4767 PAD:10471 0.0751765
rPAD/7014 PAD:4767 PAD:4770 0.0375882
rPAD/7015 PAD:4767 PAD:10475 1.5
rPAD/7016 PAD:4766 PAD:4769 0.0375882
rPAD/7017 PAD:4766 PAD:4767 1.5
rPAD/7018 PAD:4763 PAD:4766 0.0751765
rPAD/7019 PAD:4763 PAD:10471 1.5
rPAD/7020 PAD:4761 PAD:10465 0.0751765
rPAD/7021 PAD:4761 PAD:10471 0.0375882
rPAD/7022 PAD:4761 PAD:10469 1.5
rPAD/7023 PAD:4760 PAD:4763 0.0375882
rPAD/7024 PAD:4760 PAD:4761 1.5
rPAD/7025 PAD:4757 PAD:4760 0.0751765
rPAD/7026 PAD:4757 PAD:10465 1.5
rPAD/7027 PAD:4754 PAD:4757 0.0375882
rPAD/7028 PAD:4754 PAD:10462 1.5
rPAD/7029 PAD:4751 PAD:4754 0.0751765
rPAD/7030 PAD:4751 PAD:10459 1.5
rPAD/7031 PAD:4749 PAD:10453 0.0751765
rPAD/7032 PAD:4749 PAD:10459 0.0375882
rPAD/7033 PAD:4749 PAD:10457 1.5
rPAD/7034 PAD:4748 PAD:4751 0.0375882
rPAD/7035 PAD:4748 PAD:4749 1.5
rPAD/7036 PAD:4745 PAD:4748 0.0751765
rPAD/7037 PAD:4745 PAD:10453 1.5
rPAD/7038 PAD:4742 PAD:4745 0.0375882
rPAD/7039 PAD:4742 PAD:10450 1.5
rPAD/7040 PAD:4740 PAD:10450 0.0751765
rPAD/7041 PAD:4740 PAD:10448 1.5
rPAD/7042 PAD:4739 PAD:4742 0.0751765
rPAD/7043 PAD:4739 PAD:4740 1.5
rPAD/7044 PAD:4737 PAD:4740 0.0375882
rPAD/7045 PAD:4737 PAD:10445 1.5
rPAD/7046 PAD:4736 PAD:4739 0.0375882
rPAD/7047 PAD:4736 PAD:4737 1.5
rPAD/7048 PAD:4734 PAD:4737 0.0751765
rPAD/7049 PAD:4734 PAD:10442 1.5
rPAD/7050 PAD:4733 PAD:4736 0.0751765
rPAD/7051 PAD:4733 PAD:4734 1.5
rPAD/7052 PAD:4731 PAD:4734 0.0375882
rPAD/7053 PAD:4731 PAD:10439 1.5
rPAD/7054 PAD:4730 PAD:4733 0.0375882
rPAD/7055 PAD:4730 PAD:4731 1.5
rPAD/7056 PAD:4728 PAD:4731 0.0751765
rPAD/7057 PAD:4728 PAD:10436 1.5
rPAD/7058 PAD:4727 PAD:4730 0.0751765
rPAD/7059 PAD:4727 PAD:4728 1.5
rPAD/7060 PAD:4725 PAD:10429 0.0751765
rPAD/7061 PAD:4725 PAD:4728 0.0375882
rPAD/7062 PAD:4725 PAD:10433 1.5
rPAD/7063 PAD:4724 PAD:4727 0.0375882
rPAD/7064 PAD:4724 PAD:4725 1.5
rPAD/7065 PAD:4721 PAD:4724 0.0751765
rPAD/7066 PAD:4721 PAD:10429 1.5
rPAD/7067 PAD:4719 PAD:10429 0.0375882
rPAD/7068 PAD:4719 PAD:10427 1.5
rPAD/7069 PAD:4718 PAD:4721 0.0375882
rPAD/7070 PAD:4718 PAD:4719 1.5
rPAD/7071 PAD:4716 PAD:4719 0.0751765
rPAD/7072 PAD:4716 PAD:10424 1.5
rPAD/7073 PAD:4715 PAD:4718 0.0751765
rPAD/7074 PAD:4715 PAD:4716 1.5
rPAD/7075 PAD:4713 PAD:10417 0.0751765
rPAD/7076 PAD:4713 PAD:4716 0.0375882
rPAD/7077 PAD:4713 PAD:10421 1.5
rPAD/7078 PAD:4712 PAD:4715 0.0375882
rPAD/7079 PAD:4712 PAD:4713 1.5
rPAD/7080 PAD:4709 PAD:4712 0.0751765
rPAD/7081 PAD:4709 PAD:10417 1.5
rPAD/7082 PAD:4706 PAD:4709 0.0375882
rPAD/7083 PAD:4706 PAD:10414 1.5
rPAD/7084 PAD:4703 PAD:4706 0.0751765
rPAD/7085 PAD:4703 PAD:10411 1.5
rPAD/7086 PAD:4700 PAD:4703 0.0375882
rPAD/7087 PAD:4700 PAD:10408 1.5
rPAD/7088 PAD:4697 PAD:4700 0.0751765
rPAD/7089 PAD:4697 PAD:10405 1.5
rPAD/7090 PAD:4695 PAD:10405 0.0375882
rPAD/7091 PAD:4695 PAD:10403 1.5
rPAD/7092 PAD:4694 PAD:4697 0.0375882
rPAD/7093 PAD:4694 PAD:4695 1.5
rPAD/7094 PAD:4692 PAD:10396 0.0375882
rPAD/7095 PAD:4692 PAD:4695 0.0751765
rPAD/7096 PAD:4692 PAD:10400 1.5
rPAD/7097 PAD:4691 PAD:4694 0.0751765
rPAD/7098 PAD:4691 PAD:4692 1.5
rPAD/7099 PAD:4688 PAD:4691 0.0375882
rPAD/7100 PAD:4688 PAD:10396 1.5
rPAD/7101 PAD:4686 PAD:10396 0.0751765
rPAD/7102 PAD:4686 PAD:10394 1.5
rPAD/7103 PAD:4685 PAD:4688 0.0751765
rPAD/7104 PAD:4685 PAD:4686 1.5
rPAD/7105 PAD:4683 PAD:4686 0.0375882
rPAD/7106 PAD:4683 PAD:10391 1.5
rPAD/7107 PAD:4682 PAD:4685 0.0375882
rPAD/7108 PAD:4682 PAD:4683 1.5
rPAD/7109 PAD:4680 PAD:4683 0.0751765
rPAD/7110 PAD:4680 PAD:10388 1.5
rPAD/7111 PAD:4679 PAD:4682 0.0751765
rPAD/7112 PAD:4679 PAD:4680 1.5
rPAD/7113 PAD:4677 PAD:4680 0.0375882
rPAD/7114 PAD:4677 PAD:10385 1.5
rPAD/7115 PAD:4676 PAD:4679 0.0375882
rPAD/7116 PAD:4676 PAD:4677 1.5
rPAD/7117 PAD:4674 PAD:4677 0.0751765
rPAD/7118 PAD:4674 PAD:10382 1.5
rPAD/7119 PAD:4673 PAD:4676 0.0751765
rPAD/7120 PAD:4673 PAD:4674 1.5
rPAD/7121 PAD:4671 PAD:10375 0.0751765
rPAD/7122 PAD:4671 PAD:4674 0.0375882
rPAD/7123 PAD:4671 PAD:10379 1.5
rPAD/7124 PAD:4670 PAD:4673 0.0375882
rPAD/7125 PAD:4670 PAD:4671 1.5
rPAD/7126 PAD:4667 PAD:4670 0.0751765
rPAD/7127 PAD:4667 PAD:10375 1.5
rPAD/7128 PAD:4665 PAD:10375 0.0375882
rPAD/7129 PAD:4665 PAD:10373 1.5
rPAD/7130 PAD:4664 PAD:4667 0.0375882
rPAD/7131 PAD:4664 PAD:4665 1.5
rPAD/7132 PAD:4662 PAD:4665 0.0751765
rPAD/7133 PAD:4662 PAD:10370 1.5
rPAD/7134 PAD:4661 PAD:4664 0.0751765
rPAD/7135 PAD:4661 PAD:4662 1.5
rPAD/7136 PAD:4659 PAD:4662 0.0375882
rPAD/7137 PAD:4659 PAD:10367 1.5
rPAD/7138 PAD:4658 PAD:4661 0.0375882
rPAD/7139 PAD:4658 PAD:4659 1.5
rPAD/7140 PAD:4656 PAD:4659 0.0751765
rPAD/7141 PAD:4656 PAD:10364 1.5
rPAD/7142 PAD:4655 PAD:4658 0.0751765
rPAD/7143 PAD:4655 PAD:4656 1.5
rPAD/7144 PAD:4653 PAD:4656 0.0375882
rPAD/7145 PAD:4653 PAD:10361 1.5
rPAD/7146 PAD:4652 PAD:4655 0.0375882
rPAD/7147 PAD:4652 PAD:4653 1.5
rPAD/7148 PAD:4650 PAD:4653 0.0751765
rPAD/7149 PAD:4650 PAD:10358 1.5
rPAD/7150 PAD:4649 PAD:4652 0.0751765
rPAD/7151 PAD:4649 PAD:4650 1.5
rPAD/7152 PAD:4647 PAD:4650 0.0375882
rPAD/7153 PAD:4647 PAD:10355 1.5
rPAD/7154 PAD:4646 PAD:4649 0.0375882
rPAD/7155 PAD:4646 PAD:4647 1.5
rPAD/7156 PAD:4644 PAD:14857 0.0283817
rPAD/7157 PAD:4644 PAD:4647 0.0751765
rPAD/7158 PAD:4644 PAD:10352 1.5
rPAD/7159 PAD:4643 PAD:9132 0.0378785
rPAD/7160 PAD:4643 PAD:4646 0.0751765
rPAD/7161 PAD:4643 PAD:4644 1.5
rPAD/7162 PAD:4639 PAD:10179 0.0100588
rPAD/7163 PAD:4639 PAD:10347 1.5
rPAD/7164 PAD:4638 PAD:9331 0.0670908
rPAD/7165 PAD:4638 PAD:4639 1.5
rPAD/7166 PAD:4636 PAD:4639 0.0751765
rPAD/7167 PAD:4636 PAD:10344 1.5
rPAD/7168 PAD:4635 PAD:4638 0.0751765
rPAD/7169 PAD:4635 PAD:4636 1.5
rPAD/7170 PAD:4633 PAD:10337 0.0751765
rPAD/7171 PAD:4633 PAD:4636 0.0375882
rPAD/7172 PAD:4633 PAD:10341 1.5
rPAD/7173 PAD:4632 PAD:4635 0.0375882
rPAD/7174 PAD:4632 PAD:4633 1.5
rPAD/7175 PAD:4629 PAD:4632 0.0751765
rPAD/7176 PAD:4629 PAD:10337 1.5
rPAD/7177 PAD:4627 PAD:10337 0.0375882
rPAD/7178 PAD:4627 PAD:10335 1.5
rPAD/7179 PAD:4626 PAD:4629 0.0375882
rPAD/7180 PAD:4626 PAD:4627 1.5
rPAD/7181 PAD:4624 PAD:4627 0.0751765
rPAD/7182 PAD:4624 PAD:10332 1.5
rPAD/7183 PAD:4623 PAD:4626 0.0751765
rPAD/7184 PAD:4623 PAD:4624 1.5
rPAD/7185 PAD:4621 PAD:4624 0.0375882
rPAD/7186 PAD:4621 PAD:10329 1.5
rPAD/7187 PAD:4620 PAD:4623 0.0375882
rPAD/7188 PAD:4620 PAD:4621 1.5
rPAD/7189 PAD:4618 PAD:4621 0.0751765
rPAD/7190 PAD:4618 PAD:10326 1.5
rPAD/7191 PAD:4617 PAD:4620 0.0751765
rPAD/7192 PAD:4617 PAD:4618 1.5
rPAD/7193 PAD:4615 PAD:4618 0.0375882
rPAD/7194 PAD:4615 PAD:10323 1.5
rPAD/7195 PAD:4614 PAD:4617 0.0375882
rPAD/7196 PAD:4614 PAD:4615 1.5
rPAD/7197 PAD:4612 PAD:4615 0.0751765
rPAD/7198 PAD:4612 PAD:10320 1.5
rPAD/7199 PAD:4611 PAD:4614 0.0751765
rPAD/7200 PAD:4611 PAD:4612 1.5
rPAD/7201 PAD:4609 PAD:4612 0.0375882
rPAD/7202 PAD:4609 PAD:10317 1.5
rPAD/7203 PAD:4608 PAD:4611 0.0375882
rPAD/7204 PAD:4608 PAD:4609 1.5
rPAD/7205 PAD:4606 PAD:4609 0.0751765
rPAD/7206 PAD:4606 PAD:10314 1.5
rPAD/7207 PAD:4605 PAD:4608 0.0751765
rPAD/7208 PAD:4605 PAD:4606 1.5
rPAD/7209 PAD:4603 PAD:4606 0.0375882
rPAD/7210 PAD:4603 PAD:10311 1.5
rPAD/7211 PAD:4602 PAD:4605 0.0375882
rPAD/7212 PAD:4602 PAD:4603 1.5
rPAD/7213 PAD:4600 PAD:4603 0.0751765
rPAD/7214 PAD:4600 PAD:10308 1.5
rPAD/7215 PAD:4599 PAD:4602 0.0751765
rPAD/7216 PAD:4599 PAD:4600 1.5
rPAD/7217 PAD:4597 PAD:10301 0.0751765
rPAD/7218 PAD:4597 PAD:4600 0.0375882
rPAD/7219 PAD:4597 PAD:10305 1.5
rPAD/7220 PAD:4596 PAD:4599 0.0375882
rPAD/7221 PAD:4596 PAD:4597 1.5
rPAD/7222 PAD:4593 PAD:4596 0.0751765
rPAD/7223 PAD:4593 PAD:10301 1.5
rPAD/7224 PAD:4591 PAD:10295 0.0751765
rPAD/7225 PAD:4591 PAD:10301 0.0375882
rPAD/7226 PAD:4591 PAD:10299 1.5
rPAD/7227 PAD:4590 PAD:4593 0.0375882
rPAD/7228 PAD:4590 PAD:4591 1.5
rPAD/7229 PAD:4587 PAD:4590 0.0751765
rPAD/7230 PAD:4587 PAD:10295 1.5
rPAD/7231 PAD:4584 PAD:4587 0.0375882
rPAD/7232 PAD:4584 PAD:10292 1.5
rPAD/7233 PAD:4581 PAD:4584 0.0751765
rPAD/7234 PAD:4581 PAD:10289 1.5
rPAD/7235 PAD:4579 PAD:10283 0.0751765
rPAD/7236 PAD:4579 PAD:10289 0.0375882
rPAD/7237 PAD:4579 PAD:10287 1.5
rPAD/7238 PAD:4578 PAD:4581 0.0375882
rPAD/7239 PAD:4578 PAD:4579 1.5
rPAD/7240 PAD:4575 PAD:4578 0.0751765
rPAD/7241 PAD:4575 PAD:10283 1.5
rPAD/7242 PAD:4572 PAD:4575 0.0375882
rPAD/7243 PAD:4572 PAD:10280 1.5
rPAD/7244 PAD:4570 PAD:10280 0.0751765
rPAD/7245 PAD:4570 PAD:10278 1.5
rPAD/7246 PAD:4569 PAD:4572 0.0751765
rPAD/7247 PAD:4569 PAD:4570 1.5
rPAD/7248 PAD:4567 PAD:4570 0.0375882
rPAD/7249 PAD:4567 PAD:10275 1.5
rPAD/7250 PAD:4566 PAD:4569 0.0375882
rPAD/7251 PAD:4566 PAD:4567 1.5
rPAD/7252 PAD:4564 PAD:4567 0.0751765
rPAD/7253 PAD:4564 PAD:10272 1.5
rPAD/7254 PAD:4563 PAD:4566 0.0751765
rPAD/7255 PAD:4563 PAD:4564 1.5
rPAD/7256 PAD:4561 PAD:4564 0.0375882
rPAD/7257 PAD:4561 PAD:10269 1.5
rPAD/7258 PAD:4560 PAD:4563 0.0375882
rPAD/7259 PAD:4560 PAD:4561 1.5
rPAD/7260 PAD:4558 PAD:4561 0.0751765
rPAD/7261 PAD:4558 PAD:10266 1.5
rPAD/7262 PAD:4557 PAD:4560 0.0751765
rPAD/7263 PAD:4557 PAD:4558 1.5
rPAD/7264 PAD:4555 PAD:10259 0.0751765
rPAD/7265 PAD:4555 PAD:4558 0.0375882
rPAD/7266 PAD:4555 PAD:10263 1.5
rPAD/7267 PAD:4554 PAD:4557 0.0375882
rPAD/7268 PAD:4554 PAD:4555 1.5
rPAD/7269 PAD:4551 PAD:4554 0.0751765
rPAD/7270 PAD:4551 PAD:10259 1.5
rPAD/7271 PAD:4549 PAD:10259 0.0375882
rPAD/7272 PAD:4549 PAD:10257 1.5
rPAD/7273 PAD:4548 PAD:4551 0.0375882
rPAD/7274 PAD:4548 PAD:4549 1.5
rPAD/7275 PAD:4546 PAD:4549 0.0751765
rPAD/7276 PAD:4546 PAD:10254 1.5
rPAD/7277 PAD:4545 PAD:4548 0.0751765
rPAD/7278 PAD:4545 PAD:4546 1.5
rPAD/7279 PAD:4543 PAD:10247 0.0751765
rPAD/7280 PAD:4543 PAD:4546 0.0375882
rPAD/7281 PAD:4543 PAD:10251 1.5
rPAD/7282 PAD:4542 PAD:4545 0.0375882
rPAD/7283 PAD:4542 PAD:4543 1.5
rPAD/7284 PAD:4539 PAD:4542 0.0751765
rPAD/7285 PAD:4539 PAD:10247 1.5
rPAD/7286 PAD:4536 PAD:4539 0.0375882
rPAD/7287 PAD:4536 PAD:10244 1.5
rPAD/7288 PAD:4533 PAD:4536 0.0751765
rPAD/7289 PAD:4533 PAD:10241 1.5
rPAD/7290 PAD:4530 PAD:4533 0.0375882
rPAD/7291 PAD:4530 PAD:10238 1.5
rPAD/7292 PAD:4527 PAD:4530 0.0751765
rPAD/7293 PAD:4527 PAD:10235 1.5
rPAD/7294 PAD:4525 PAD:10235 0.0375882
rPAD/7295 PAD:4525 PAD:10233 1.5
rPAD/7296 PAD:4524 PAD:4527 0.0375882
rPAD/7297 PAD:4524 PAD:4525 1.5
rPAD/7298 PAD:4522 PAD:10226 0.0375882
rPAD/7299 PAD:4522 PAD:4525 0.0751765
rPAD/7300 PAD:4522 PAD:10230 1.5
rPAD/7301 PAD:4521 PAD:4524 0.0751765
rPAD/7302 PAD:4521 PAD:4522 1.5
rPAD/7303 PAD:4518 PAD:4521 0.0375882
rPAD/7304 PAD:4518 PAD:10226 1.5
rPAD/7305 PAD:4516 PAD:10226 0.0751765
rPAD/7306 PAD:4516 PAD:10224 1.5
rPAD/7307 PAD:4515 PAD:4518 0.0751765
rPAD/7308 PAD:4515 PAD:4516 1.5
rPAD/7309 PAD:4513 PAD:4516 0.0375882
rPAD/7310 PAD:4513 PAD:10221 1.5
rPAD/7311 PAD:4512 PAD:4515 0.0375882
rPAD/7312 PAD:4512 PAD:4513 1.5
rPAD/7313 PAD:4510 PAD:4513 0.0751765
rPAD/7314 PAD:4510 PAD:10218 1.5
rPAD/7315 PAD:4509 PAD:4512 0.0751765
rPAD/7316 PAD:4509 PAD:4510 1.5
rPAD/7317 PAD:4507 PAD:4510 0.0375882
rPAD/7318 PAD:4507 PAD:10215 1.5
rPAD/7319 PAD:4506 PAD:4509 0.0375882
rPAD/7320 PAD:4506 PAD:4507 1.5
rPAD/7321 PAD:4504 PAD:4507 0.0751765
rPAD/7322 PAD:4504 PAD:10212 1.5
rPAD/7323 PAD:4503 PAD:4506 0.0751765
rPAD/7324 PAD:4503 PAD:4504 1.5
rPAD/7325 PAD:4501 PAD:10205 0.0751765
rPAD/7326 PAD:4501 PAD:4504 0.0375882
rPAD/7327 PAD:4501 PAD:10209 1.5
rPAD/7328 PAD:4500 PAD:4503 0.0375882
rPAD/7329 PAD:4500 PAD:4501 1.5
rPAD/7330 PAD:4497 PAD:4500 0.0751765
rPAD/7331 PAD:4497 PAD:10205 1.5
rPAD/7332 PAD:4495 PAD:10205 0.0375882
rPAD/7333 PAD:4495 PAD:10203 1.5
rPAD/7334 PAD:4494 PAD:4497 0.0375882
rPAD/7335 PAD:4494 PAD:4495 1.5
rPAD/7336 PAD:4492 PAD:4495 0.0751765
rPAD/7337 PAD:4492 PAD:10200 1.5
rPAD/7338 PAD:4491 PAD:4494 0.0751765
rPAD/7339 PAD:4491 PAD:4492 1.5
rPAD/7340 PAD:4489 PAD:4492 0.0375882
rPAD/7341 PAD:4489 PAD:10197 1.5
rPAD/7342 PAD:4488 PAD:4491 0.0375882
rPAD/7343 PAD:4488 PAD:4489 1.5
rPAD/7344 PAD:4486 PAD:4489 0.0751765
rPAD/7345 PAD:4486 PAD:10194 1.5
rPAD/7346 PAD:4485 PAD:4488 0.0751765
rPAD/7347 PAD:4485 PAD:4486 1.5
rPAD/7348 PAD:4483 PAD:4486 0.0375882
rPAD/7349 PAD:4483 PAD:10191 1.5
rPAD/7350 PAD:4482 PAD:4485 0.0375882
rPAD/7351 PAD:4482 PAD:4483 1.5
rPAD/7352 PAD:4480 PAD:4483 0.0751765
rPAD/7353 PAD:4480 PAD:10188 1.5
rPAD/7354 PAD:4479 PAD:4482 0.0751765
rPAD/7355 PAD:4479 PAD:4480 1.5
rPAD/7356 PAD:4477 PAD:4480 0.0375882
rPAD/7357 PAD:4477 PAD:10185 1.5
rPAD/7358 PAD:4476 PAD:4479 0.0375882
rPAD/7359 PAD:4476 PAD:4477 1.5
rPAD/7360 PAD:4474 PAD:14852 0.0283817
rPAD/7361 PAD:4474 PAD:4477 0.0751765
rPAD/7362 PAD:4474 PAD:10182 1.5
rPAD/7363 PAD:4473 PAD:9125 0.0378785
rPAD/7364 PAD:4473 PAD:4476 0.0751765
rPAD/7365 PAD:4473 PAD:4474 1.5
rPAD/7366 PAD:4469 PAD:10009 0.0100588
rPAD/7367 PAD:4469 PAD:10177 1.5
rPAD/7368 PAD:4468 PAD:9327 0.0670908
rPAD/7369 PAD:4468 PAD:4469 1.5
rPAD/7370 PAD:4466 PAD:4469 0.0751765
rPAD/7371 PAD:4466 PAD:10174 1.5
rPAD/7372 PAD:4465 PAD:4468 0.0751765
rPAD/7373 PAD:4465 PAD:4466 1.5
rPAD/7374 PAD:4463 PAD:10167 0.0751765
rPAD/7375 PAD:4463 PAD:4466 0.0375882
rPAD/7376 PAD:4463 PAD:10171 1.5
rPAD/7377 PAD:4462 PAD:4465 0.0375882
rPAD/7378 PAD:4462 PAD:4463 1.5
rPAD/7379 PAD:4459 PAD:4462 0.0751765
rPAD/7380 PAD:4459 PAD:10167 1.5
rPAD/7381 PAD:4457 PAD:10167 0.0375882
rPAD/7382 PAD:4457 PAD:10165 1.5
rPAD/7383 PAD:4456 PAD:4459 0.0375882
rPAD/7384 PAD:4456 PAD:4457 1.5
rPAD/7385 PAD:4454 PAD:4457 0.0751765
rPAD/7386 PAD:4454 PAD:10162 1.5
rPAD/7387 PAD:4453 PAD:4456 0.0751765
rPAD/7388 PAD:4453 PAD:4454 1.5
rPAD/7389 PAD:4451 PAD:4454 0.0375882
rPAD/7390 PAD:4451 PAD:10159 1.5
rPAD/7391 PAD:4450 PAD:4453 0.0375882
rPAD/7392 PAD:4450 PAD:4451 1.5
rPAD/7393 PAD:4448 PAD:4451 0.0751765
rPAD/7394 PAD:4448 PAD:10156 1.5
rPAD/7395 PAD:4447 PAD:4450 0.0751765
rPAD/7396 PAD:4447 PAD:4448 1.5
rPAD/7397 PAD:4445 PAD:4448 0.0375882
rPAD/7398 PAD:4445 PAD:10153 1.5
rPAD/7399 PAD:4444 PAD:4447 0.0375882
rPAD/7400 PAD:4444 PAD:4445 1.5
rPAD/7401 PAD:4442 PAD:4445 0.0751765
rPAD/7402 PAD:4442 PAD:10150 1.5
rPAD/7403 PAD:4441 PAD:4444 0.0751765
rPAD/7404 PAD:4441 PAD:4442 1.5
rPAD/7405 PAD:4439 PAD:4442 0.0375882
rPAD/7406 PAD:4439 PAD:10147 1.5
rPAD/7407 PAD:4438 PAD:4441 0.0375882
rPAD/7408 PAD:4438 PAD:4439 1.5
rPAD/7409 PAD:4436 PAD:4439 0.0751765
rPAD/7410 PAD:4436 PAD:10144 1.5
rPAD/7411 PAD:4435 PAD:4438 0.0751765
rPAD/7412 PAD:4435 PAD:4436 1.5
rPAD/7413 PAD:4433 PAD:4436 0.0375882
rPAD/7414 PAD:4433 PAD:10141 1.5
rPAD/7415 PAD:4432 PAD:4435 0.0375882
rPAD/7416 PAD:4432 PAD:4433 1.5
rPAD/7417 PAD:4430 PAD:4433 0.0751765
rPAD/7418 PAD:4430 PAD:10138 1.5
rPAD/7419 PAD:4429 PAD:4432 0.0751765
rPAD/7420 PAD:4429 PAD:4430 1.5
rPAD/7421 PAD:4427 PAD:10131 0.0751765
rPAD/7422 PAD:4427 PAD:4430 0.0375882
rPAD/7423 PAD:4427 PAD:10135 1.5
rPAD/7424 PAD:4426 PAD:4429 0.0375882
rPAD/7425 PAD:4426 PAD:4427 1.5
rPAD/7426 PAD:4423 PAD:4426 0.0751765
rPAD/7427 PAD:4423 PAD:10131 1.5
rPAD/7428 PAD:4421 PAD:10125 0.0751765
rPAD/7429 PAD:4421 PAD:10131 0.0375882
rPAD/7430 PAD:4421 PAD:10129 1.5
rPAD/7431 PAD:4420 PAD:4423 0.0375882
rPAD/7432 PAD:4420 PAD:4421 1.5
rPAD/7433 PAD:4417 PAD:4420 0.0751765
rPAD/7434 PAD:4417 PAD:10125 1.5
rPAD/7435 PAD:4414 PAD:4417 0.0375882
rPAD/7436 PAD:4414 PAD:10122 1.5
rPAD/7437 PAD:4411 PAD:4414 0.0751765
rPAD/7438 PAD:4411 PAD:10119 1.5
rPAD/7439 PAD:4409 PAD:10113 0.0751765
rPAD/7440 PAD:4409 PAD:10119 0.0375882
rPAD/7441 PAD:4409 PAD:10117 1.5
rPAD/7442 PAD:4408 PAD:4411 0.0375882
rPAD/7443 PAD:4408 PAD:4409 1.5
rPAD/7444 PAD:4405 PAD:4408 0.0751765
rPAD/7445 PAD:4405 PAD:10113 1.5
rPAD/7446 PAD:4402 PAD:4405 0.0375882
rPAD/7447 PAD:4402 PAD:10110 1.5
rPAD/7448 PAD:4400 PAD:10110 0.0751765
rPAD/7449 PAD:4400 PAD:10108 1.5
rPAD/7450 PAD:4399 PAD:4402 0.0751765
rPAD/7451 PAD:4399 PAD:4400 1.5
rPAD/7452 PAD:4397 PAD:4400 0.0375882
rPAD/7453 PAD:4397 PAD:10105 1.5
rPAD/7454 PAD:4396 PAD:4399 0.0375882
rPAD/7455 PAD:4396 PAD:4397 1.5
rPAD/7456 PAD:4394 PAD:4397 0.0751765
rPAD/7457 PAD:4394 PAD:10102 1.5
rPAD/7458 PAD:4393 PAD:4396 0.0751765
rPAD/7459 PAD:4393 PAD:4394 1.5
rPAD/7460 PAD:4391 PAD:4394 0.0375882
rPAD/7461 PAD:4391 PAD:10099 1.5
rPAD/7462 PAD:4390 PAD:4393 0.0375882
rPAD/7463 PAD:4390 PAD:4391 1.5
rPAD/7464 PAD:4388 PAD:4391 0.0751765
rPAD/7465 PAD:4388 PAD:10096 1.5
rPAD/7466 PAD:4387 PAD:4390 0.0751765
rPAD/7467 PAD:4387 PAD:4388 1.5
rPAD/7468 PAD:4385 PAD:10089 0.0751765
rPAD/7469 PAD:4385 PAD:4388 0.0375882
rPAD/7470 PAD:4385 PAD:10093 1.5
rPAD/7471 PAD:4384 PAD:4387 0.0375882
rPAD/7472 PAD:4384 PAD:4385 1.5
rPAD/7473 PAD:4381 PAD:4384 0.0751765
rPAD/7474 PAD:4381 PAD:10089 1.5
rPAD/7475 PAD:4379 PAD:10089 0.0375882
rPAD/7476 PAD:4379 PAD:10087 1.5
rPAD/7477 PAD:4378 PAD:4381 0.0375882
rPAD/7478 PAD:4378 PAD:4379 1.5
rPAD/7479 PAD:4376 PAD:4379 0.0751765
rPAD/7480 PAD:4376 PAD:10084 1.5
rPAD/7481 PAD:4375 PAD:4378 0.0751765
rPAD/7482 PAD:4375 PAD:4376 1.5
rPAD/7483 PAD:4373 PAD:10077 0.0751765
rPAD/7484 PAD:4373 PAD:4376 0.0375882
rPAD/7485 PAD:4373 PAD:10081 1.5
rPAD/7486 PAD:4372 PAD:4375 0.0375882
rPAD/7487 PAD:4372 PAD:4373 1.5
rPAD/7488 PAD:4369 PAD:4372 0.0751765
rPAD/7489 PAD:4369 PAD:10077 1.5
rPAD/7490 PAD:4366 PAD:4369 0.0375882
rPAD/7491 PAD:4366 PAD:10074 1.5
rPAD/7492 PAD:4363 PAD:4366 0.0751765
rPAD/7493 PAD:4363 PAD:10071 1.5
rPAD/7494 PAD:4360 PAD:4363 0.0375882
rPAD/7495 PAD:4360 PAD:10068 1.5
rPAD/7496 PAD:4357 PAD:4360 0.0751765
rPAD/7497 PAD:4357 PAD:10065 1.5
rPAD/7498 PAD:4355 PAD:10065 0.0375882
rPAD/7499 PAD:4355 PAD:10063 1.5
rPAD/7500 PAD:4354 PAD:4357 0.0375882
rPAD/7501 PAD:4354 PAD:4355 1.5
rPAD/7502 PAD:4352 PAD:10056 0.0375882
rPAD/7503 PAD:4352 PAD:4355 0.0751765
rPAD/7504 PAD:4352 PAD:10060 1.5
rPAD/7505 PAD:4351 PAD:4354 0.0751765
rPAD/7506 PAD:4351 PAD:4352 1.5
rPAD/7507 PAD:4348 PAD:4351 0.0375882
rPAD/7508 PAD:4348 PAD:10056 1.5
rPAD/7509 PAD:4346 PAD:10056 0.0751765
rPAD/7510 PAD:4346 PAD:10054 1.5
rPAD/7511 PAD:4345 PAD:4348 0.0751765
rPAD/7512 PAD:4345 PAD:4346 1.5
rPAD/7513 PAD:4343 PAD:4346 0.0375882
rPAD/7514 PAD:4343 PAD:10051 1.5
rPAD/7515 PAD:4342 PAD:4345 0.0375882
rPAD/7516 PAD:4342 PAD:4343 1.5
rPAD/7517 PAD:4340 PAD:4343 0.0751765
rPAD/7518 PAD:4340 PAD:10048 1.5
rPAD/7519 PAD:4339 PAD:4342 0.0751765
rPAD/7520 PAD:4339 PAD:4340 1.5
rPAD/7521 PAD:4337 PAD:4340 0.0375882
rPAD/7522 PAD:4337 PAD:10045 1.5
rPAD/7523 PAD:4336 PAD:4339 0.0375882
rPAD/7524 PAD:4336 PAD:4337 1.5
rPAD/7525 PAD:4334 PAD:4337 0.0751765
rPAD/7526 PAD:4334 PAD:10042 1.5
rPAD/7527 PAD:4333 PAD:4336 0.0751765
rPAD/7528 PAD:4333 PAD:4334 1.5
rPAD/7529 PAD:4331 PAD:10035 0.0751765
rPAD/7530 PAD:4331 PAD:4334 0.0375882
rPAD/7531 PAD:4331 PAD:10039 1.5
rPAD/7532 PAD:4330 PAD:4333 0.0375882
rPAD/7533 PAD:4330 PAD:4331 1.5
rPAD/7534 PAD:4327 PAD:4330 0.0751765
rPAD/7535 PAD:4327 PAD:10035 1.5
rPAD/7536 PAD:4325 PAD:10035 0.0375882
rPAD/7537 PAD:4325 PAD:10033 1.5
rPAD/7538 PAD:4324 PAD:4327 0.0375882
rPAD/7539 PAD:4324 PAD:4325 1.5
rPAD/7540 PAD:4322 PAD:4325 0.0751765
rPAD/7541 PAD:4322 PAD:10030 1.5
rPAD/7542 PAD:4321 PAD:4324 0.0751765
rPAD/7543 PAD:4321 PAD:4322 1.5
rPAD/7544 PAD:4319 PAD:4322 0.0375882
rPAD/7545 PAD:4319 PAD:10027 1.5
rPAD/7546 PAD:4318 PAD:4321 0.0375882
rPAD/7547 PAD:4318 PAD:4319 1.5
rPAD/7548 PAD:4316 PAD:4319 0.0751765
rPAD/7549 PAD:4316 PAD:10024 1.5
rPAD/7550 PAD:4315 PAD:4318 0.0751765
rPAD/7551 PAD:4315 PAD:4316 1.5
rPAD/7552 PAD:4313 PAD:4316 0.0375882
rPAD/7553 PAD:4313 PAD:10021 1.5
rPAD/7554 PAD:4312 PAD:4315 0.0375882
rPAD/7555 PAD:4312 PAD:4313 1.5
rPAD/7556 PAD:4310 PAD:4313 0.0751765
rPAD/7557 PAD:4310 PAD:10018 1.5
rPAD/7558 PAD:4309 PAD:4312 0.0751765
rPAD/7559 PAD:4309 PAD:4310 1.5
rPAD/7560 PAD:4307 PAD:4310 0.0375882
rPAD/7561 PAD:4307 PAD:10015 1.5
rPAD/7562 PAD:4306 PAD:4309 0.0375882
rPAD/7563 PAD:4306 PAD:4307 1.5
rPAD/7564 PAD:4304 PAD:14847 0.0283817
rPAD/7565 PAD:4304 PAD:4307 0.0751765
rPAD/7566 PAD:4304 PAD:10012 1.5
rPAD/7567 PAD:4303 PAD:9118 0.0378785
rPAD/7568 PAD:4303 PAD:4306 0.0751765
rPAD/7569 PAD:4303 PAD:4304 1.5
rPAD/7570 PAD:4299 PAD:9839 0.0100588
rPAD/7571 PAD:4299 PAD:10007 1.5
rPAD/7572 PAD:4298 PAD:9323 0.0670908
rPAD/7573 PAD:4298 PAD:4299 1.5
rPAD/7574 PAD:4296 PAD:4299 0.0751765
rPAD/7575 PAD:4296 PAD:10004 1.5
rPAD/7576 PAD:4295 PAD:4298 0.0751765
rPAD/7577 PAD:4295 PAD:4296 1.5
rPAD/7578 PAD:4293 PAD:9997 0.0751765
rPAD/7579 PAD:4293 PAD:4296 0.0375882
rPAD/7580 PAD:4293 PAD:10001 1.5
rPAD/7581 PAD:4292 PAD:4295 0.0375882
rPAD/7582 PAD:4292 PAD:4293 1.5
rPAD/7583 PAD:4289 PAD:4292 0.0751765
rPAD/7584 PAD:4289 PAD:9997 1.5
rPAD/7585 PAD:4287 PAD:9997 0.0375882
rPAD/7586 PAD:4287 PAD:9995 1.5
rPAD/7587 PAD:4286 PAD:4289 0.0375882
rPAD/7588 PAD:4286 PAD:4287 1.5
rPAD/7589 PAD:4284 PAD:4287 0.0751765
rPAD/7590 PAD:4284 PAD:9992 1.5
rPAD/7591 PAD:4283 PAD:4286 0.0751765
rPAD/7592 PAD:4283 PAD:4284 1.5
rPAD/7593 PAD:4281 PAD:4284 0.0375882
rPAD/7594 PAD:4281 PAD:9989 1.5
rPAD/7595 PAD:4280 PAD:4283 0.0375882
rPAD/7596 PAD:4280 PAD:4281 1.5
rPAD/7597 PAD:4278 PAD:4281 0.0751765
rPAD/7598 PAD:4278 PAD:9986 1.5
rPAD/7599 PAD:4277 PAD:4280 0.0751765
rPAD/7600 PAD:4277 PAD:4278 1.5
rPAD/7601 PAD:4275 PAD:4278 0.0375882
rPAD/7602 PAD:4275 PAD:9983 1.5
rPAD/7603 PAD:4274 PAD:4277 0.0375882
rPAD/7604 PAD:4274 PAD:4275 1.5
rPAD/7605 PAD:4272 PAD:4275 0.0751765
rPAD/7606 PAD:4272 PAD:9980 1.5
rPAD/7607 PAD:4271 PAD:4274 0.0751765
rPAD/7608 PAD:4271 PAD:4272 1.5
rPAD/7609 PAD:4269 PAD:4272 0.0375882
rPAD/7610 PAD:4269 PAD:9977 1.5
rPAD/7611 PAD:4268 PAD:4271 0.0375882
rPAD/7612 PAD:4268 PAD:4269 1.5
rPAD/7613 PAD:4266 PAD:4269 0.0751765
rPAD/7614 PAD:4266 PAD:9974 1.5
rPAD/7615 PAD:4265 PAD:4268 0.0751765
rPAD/7616 PAD:4265 PAD:4266 1.5
rPAD/7617 PAD:4263 PAD:4266 0.0375882
rPAD/7618 PAD:4263 PAD:9971 1.5
rPAD/7619 PAD:4262 PAD:4265 0.0375882
rPAD/7620 PAD:4262 PAD:4263 1.5
rPAD/7621 PAD:4260 PAD:4263 0.0751765
rPAD/7622 PAD:4260 PAD:9968 1.5
rPAD/7623 PAD:4259 PAD:4262 0.0751765
rPAD/7624 PAD:4259 PAD:4260 1.5
rPAD/7625 PAD:4257 PAD:9961 0.0751765
rPAD/7626 PAD:4257 PAD:4260 0.0375882
rPAD/7627 PAD:4257 PAD:9965 1.5
rPAD/7628 PAD:4256 PAD:4259 0.0375882
rPAD/7629 PAD:4256 PAD:4257 1.5
rPAD/7630 PAD:4253 PAD:4256 0.0751765
rPAD/7631 PAD:4253 PAD:9961 1.5
rPAD/7632 PAD:4251 PAD:9955 0.0751765
rPAD/7633 PAD:4251 PAD:9961 0.0375882
rPAD/7634 PAD:4251 PAD:9959 1.5
rPAD/7635 PAD:4250 PAD:4253 0.0375882
rPAD/7636 PAD:4250 PAD:4251 1.5
rPAD/7637 PAD:4247 PAD:4250 0.0751765
rPAD/7638 PAD:4247 PAD:9955 1.5
rPAD/7639 PAD:4244 PAD:4247 0.0375882
rPAD/7640 PAD:4244 PAD:9952 1.5
rPAD/7641 PAD:4241 PAD:4244 0.0751765
rPAD/7642 PAD:4241 PAD:9949 1.5
rPAD/7643 PAD:4239 PAD:9943 0.0751765
rPAD/7644 PAD:4239 PAD:9949 0.0375882
rPAD/7645 PAD:4239 PAD:9947 1.5
rPAD/7646 PAD:4238 PAD:4241 0.0375882
rPAD/7647 PAD:4238 PAD:4239 1.5
rPAD/7648 PAD:4235 PAD:4238 0.0751765
rPAD/7649 PAD:4235 PAD:9943 1.5
rPAD/7650 PAD:4232 PAD:4235 0.0375882
rPAD/7651 PAD:4232 PAD:9940 1.5
rPAD/7652 PAD:4230 PAD:9940 0.0751765
rPAD/7653 PAD:4230 PAD:9938 1.5
rPAD/7654 PAD:4229 PAD:4232 0.0751765
rPAD/7655 PAD:4229 PAD:4230 1.5
rPAD/7656 PAD:4227 PAD:4230 0.0375882
rPAD/7657 PAD:4227 PAD:9935 1.5
rPAD/7658 PAD:4226 PAD:4229 0.0375882
rPAD/7659 PAD:4226 PAD:4227 1.5
rPAD/7660 PAD:4224 PAD:4227 0.0751765
rPAD/7661 PAD:4224 PAD:9932 1.5
rPAD/7662 PAD:4223 PAD:4226 0.0751765
rPAD/7663 PAD:4223 PAD:4224 1.5
rPAD/7664 PAD:4221 PAD:4224 0.0375882
rPAD/7665 PAD:4221 PAD:9929 1.5
rPAD/7666 PAD:4220 PAD:4223 0.0375882
rPAD/7667 PAD:4220 PAD:4221 1.5
rPAD/7668 PAD:4218 PAD:4221 0.0751765
rPAD/7669 PAD:4218 PAD:9926 1.5
rPAD/7670 PAD:4217 PAD:4220 0.0751765
rPAD/7671 PAD:4217 PAD:4218 1.5
rPAD/7672 PAD:4215 PAD:9919 0.0751765
rPAD/7673 PAD:4215 PAD:4218 0.0375882
rPAD/7674 PAD:4215 PAD:9923 1.5
rPAD/7675 PAD:4214 PAD:4217 0.0375882
rPAD/7676 PAD:4214 PAD:4215 1.5
rPAD/7677 PAD:4211 PAD:4214 0.0751765
rPAD/7678 PAD:4211 PAD:9919 1.5
rPAD/7679 PAD:4209 PAD:9919 0.0375882
rPAD/7680 PAD:4209 PAD:9917 1.5
rPAD/7681 PAD:4208 PAD:4211 0.0375882
rPAD/7682 PAD:4208 PAD:4209 1.5
rPAD/7683 PAD:4206 PAD:4209 0.0751765
rPAD/7684 PAD:4206 PAD:9914 1.5
rPAD/7685 PAD:4205 PAD:4208 0.0751765
rPAD/7686 PAD:4205 PAD:4206 1.5
rPAD/7687 PAD:4203 PAD:9907 0.0751765
rPAD/7688 PAD:4203 PAD:4206 0.0375882
rPAD/7689 PAD:4203 PAD:9911 1.5
rPAD/7690 PAD:4202 PAD:4205 0.0375882
rPAD/7691 PAD:4202 PAD:4203 1.5
rPAD/7692 PAD:4199 PAD:4202 0.0751765
rPAD/7693 PAD:4199 PAD:9907 1.5
rPAD/7694 PAD:4196 PAD:4199 0.0375882
rPAD/7695 PAD:4196 PAD:9904 1.5
rPAD/7696 PAD:4193 PAD:4196 0.0751765
rPAD/7697 PAD:4193 PAD:9901 1.5
rPAD/7698 PAD:4190 PAD:4193 0.0375882
rPAD/7699 PAD:4190 PAD:9898 1.5
rPAD/7700 PAD:4187 PAD:4190 0.0751765
rPAD/7701 PAD:4187 PAD:9895 1.5
rPAD/7702 PAD:4185 PAD:9895 0.0375882
rPAD/7703 PAD:4185 PAD:9893 1.5
rPAD/7704 PAD:4184 PAD:4187 0.0375882
rPAD/7705 PAD:4184 PAD:4185 1.5
rPAD/7706 PAD:4182 PAD:9886 0.0375882
rPAD/7707 PAD:4182 PAD:4185 0.0751765
rPAD/7708 PAD:4182 PAD:9890 1.5
rPAD/7709 PAD:4181 PAD:4184 0.0751765
rPAD/7710 PAD:4181 PAD:4182 1.5
rPAD/7711 PAD:4178 PAD:4181 0.0375882
rPAD/7712 PAD:4178 PAD:9886 1.5
rPAD/7713 PAD:4176 PAD:9886 0.0751765
rPAD/7714 PAD:4176 PAD:9884 1.5
rPAD/7715 PAD:4175 PAD:4178 0.0751765
rPAD/7716 PAD:4175 PAD:4176 1.5
rPAD/7717 PAD:4173 PAD:4176 0.0375882
rPAD/7718 PAD:4173 PAD:9881 1.5
rPAD/7719 PAD:4172 PAD:4175 0.0375882
rPAD/7720 PAD:4172 PAD:4173 1.5
rPAD/7721 PAD:4170 PAD:4173 0.0751765
rPAD/7722 PAD:4170 PAD:9878 1.5
rPAD/7723 PAD:4169 PAD:4172 0.0751765
rPAD/7724 PAD:4169 PAD:4170 1.5
rPAD/7725 PAD:4167 PAD:4170 0.0375882
rPAD/7726 PAD:4167 PAD:9875 1.5
rPAD/7727 PAD:4166 PAD:4169 0.0375882
rPAD/7728 PAD:4166 PAD:4167 1.5
rPAD/7729 PAD:4164 PAD:4167 0.0751765
rPAD/7730 PAD:4164 PAD:9872 1.5
rPAD/7731 PAD:4163 PAD:4166 0.0751765
rPAD/7732 PAD:4163 PAD:4164 1.5
rPAD/7733 PAD:4161 PAD:9865 0.0751765
rPAD/7734 PAD:4161 PAD:4164 0.0375882
rPAD/7735 PAD:4161 PAD:9869 1.5
rPAD/7736 PAD:4160 PAD:4163 0.0375882
rPAD/7737 PAD:4160 PAD:4161 1.5
rPAD/7738 PAD:4157 PAD:4160 0.0751765
rPAD/7739 PAD:4157 PAD:9865 1.5
rPAD/7740 PAD:4155 PAD:9865 0.0375882
rPAD/7741 PAD:4155 PAD:9863 1.5
rPAD/7742 PAD:4154 PAD:4157 0.0375882
rPAD/7743 PAD:4154 PAD:4155 1.5
rPAD/7744 PAD:4152 PAD:4155 0.0751765
rPAD/7745 PAD:4152 PAD:9860 1.5
rPAD/7746 PAD:4151 PAD:4154 0.0751765
rPAD/7747 PAD:4151 PAD:4152 1.5
rPAD/7748 PAD:4149 PAD:4152 0.0375882
rPAD/7749 PAD:4149 PAD:9857 1.5
rPAD/7750 PAD:4148 PAD:4151 0.0375882
rPAD/7751 PAD:4148 PAD:4149 1.5
rPAD/7752 PAD:4146 PAD:4149 0.0751765
rPAD/7753 PAD:4146 PAD:9854 1.5
rPAD/7754 PAD:4145 PAD:4148 0.0751765
rPAD/7755 PAD:4145 PAD:4146 1.5
rPAD/7756 PAD:4143 PAD:4146 0.0375882
rPAD/7757 PAD:4143 PAD:9851 1.5
rPAD/7758 PAD:4142 PAD:4145 0.0375882
rPAD/7759 PAD:4142 PAD:4143 1.5
rPAD/7760 PAD:4140 PAD:4143 0.0751765
rPAD/7761 PAD:4140 PAD:9848 1.5
rPAD/7762 PAD:4139 PAD:4142 0.0751765
rPAD/7763 PAD:4139 PAD:4140 1.5
rPAD/7764 PAD:4137 PAD:4140 0.0375882
rPAD/7765 PAD:4137 PAD:9845 1.5
rPAD/7766 PAD:4136 PAD:4139 0.0375882
rPAD/7767 PAD:4136 PAD:4137 1.5
rPAD/7768 PAD:4134 PAD:14839 0.0283817
rPAD/7769 PAD:4134 PAD:4137 0.0751765
rPAD/7770 PAD:4134 PAD:9842 1.5
rPAD/7771 PAD:4133 PAD:9111 0.0378785
rPAD/7772 PAD:4133 PAD:4136 0.0751765
rPAD/7773 PAD:4133 PAD:4134 1.5
rPAD/7774 PAD:4129 PAD:9669 0.0100588
rPAD/7775 PAD:4129 PAD:9837 1.5
rPAD/7776 PAD:4128 PAD:9319 0.0670908
rPAD/7777 PAD:4128 PAD:4129 1.5
rPAD/7778 PAD:4126 PAD:4129 0.0751765
rPAD/7779 PAD:4126 PAD:9834 1.5
rPAD/7780 PAD:4125 PAD:4128 0.0751765
rPAD/7781 PAD:4125 PAD:4126 1.5
rPAD/7782 PAD:4123 PAD:9827 0.0751765
rPAD/7783 PAD:4123 PAD:4126 0.0375882
rPAD/7784 PAD:4123 PAD:9831 1.5
rPAD/7785 PAD:4122 PAD:4125 0.0375882
rPAD/7786 PAD:4122 PAD:4123 1.5
rPAD/7787 PAD:4119 PAD:4122 0.0751765
rPAD/7788 PAD:4119 PAD:9827 1.5
rPAD/7789 PAD:4117 PAD:9827 0.0375882
rPAD/7790 PAD:4117 PAD:9825 1.5
rPAD/7791 PAD:4116 PAD:4119 0.0375882
rPAD/7792 PAD:4116 PAD:4117 1.5
rPAD/7793 PAD:4114 PAD:4117 0.0751765
rPAD/7794 PAD:4114 PAD:9822 1.5
rPAD/7795 PAD:4113 PAD:4116 0.0751765
rPAD/7796 PAD:4113 PAD:4114 1.5
rPAD/7797 PAD:4111 PAD:4114 0.0375882
rPAD/7798 PAD:4111 PAD:9819 1.5
rPAD/7799 PAD:4110 PAD:4113 0.0375882
rPAD/7800 PAD:4110 PAD:4111 1.5
rPAD/7801 PAD:4108 PAD:4111 0.0751765
rPAD/7802 PAD:4108 PAD:9816 1.5
rPAD/7803 PAD:4107 PAD:4110 0.0751765
rPAD/7804 PAD:4107 PAD:4108 1.5
rPAD/7805 PAD:4105 PAD:4108 0.0375882
rPAD/7806 PAD:4105 PAD:9813 1.5
rPAD/7807 PAD:4104 PAD:4107 0.0375882
rPAD/7808 PAD:4104 PAD:4105 1.5
rPAD/7809 PAD:4102 PAD:4105 0.0751765
rPAD/7810 PAD:4102 PAD:9810 1.5
rPAD/7811 PAD:4101 PAD:4104 0.0751765
rPAD/7812 PAD:4101 PAD:4102 1.5
rPAD/7813 PAD:4099 PAD:4102 0.0375882
rPAD/7814 PAD:4099 PAD:9807 1.5
rPAD/7815 PAD:4098 PAD:4101 0.0375882
rPAD/7816 PAD:4098 PAD:4099 1.5
rPAD/7817 PAD:4096 PAD:4099 0.0751765
rPAD/7818 PAD:4096 PAD:9804 1.5
rPAD/7819 PAD:4095 PAD:4098 0.0751765
rPAD/7820 PAD:4095 PAD:4096 1.5
rPAD/7821 PAD:4093 PAD:4096 0.0375882
rPAD/7822 PAD:4093 PAD:9801 1.5
rPAD/7823 PAD:4092 PAD:4095 0.0375882
rPAD/7824 PAD:4092 PAD:4093 1.5
rPAD/7825 PAD:4090 PAD:4093 0.0751765
rPAD/7826 PAD:4090 PAD:9798 1.5
rPAD/7827 PAD:4089 PAD:4092 0.0751765
rPAD/7828 PAD:4089 PAD:4090 1.5
rPAD/7829 PAD:4087 PAD:9791 0.0751765
rPAD/7830 PAD:4087 PAD:4090 0.0375882
rPAD/7831 PAD:4087 PAD:9795 1.5
rPAD/7832 PAD:4086 PAD:4089 0.0375882
rPAD/7833 PAD:4086 PAD:4087 1.5
rPAD/7834 PAD:4083 PAD:4086 0.0751765
rPAD/7835 PAD:4083 PAD:9791 1.5
rPAD/7836 PAD:4081 PAD:9785 0.0751765
rPAD/7837 PAD:4081 PAD:9791 0.0375882
rPAD/7838 PAD:4081 PAD:9789 1.5
rPAD/7839 PAD:4080 PAD:4083 0.0375882
rPAD/7840 PAD:4080 PAD:4081 1.5
rPAD/7841 PAD:4077 PAD:4080 0.0751765
rPAD/7842 PAD:4077 PAD:9785 1.5
rPAD/7843 PAD:4074 PAD:4077 0.0375882
rPAD/7844 PAD:4074 PAD:9782 1.5
rPAD/7845 PAD:4071 PAD:4074 0.0751765
rPAD/7846 PAD:4071 PAD:9779 1.5
rPAD/7847 PAD:4069 PAD:9773 0.0751765
rPAD/7848 PAD:4069 PAD:9779 0.0375882
rPAD/7849 PAD:4069 PAD:9777 1.5
rPAD/7850 PAD:4068 PAD:4071 0.0375882
rPAD/7851 PAD:4068 PAD:4069 1.5
rPAD/7852 PAD:4065 PAD:4068 0.0751765
rPAD/7853 PAD:4065 PAD:9773 1.5
rPAD/7854 PAD:4062 PAD:4065 0.0375882
rPAD/7855 PAD:4062 PAD:9770 1.5
rPAD/7856 PAD:4060 PAD:9770 0.0751765
rPAD/7857 PAD:4060 PAD:9768 1.5
rPAD/7858 PAD:4059 PAD:4062 0.0751765
rPAD/7859 PAD:4059 PAD:4060 1.5
rPAD/7860 PAD:4057 PAD:4060 0.0375882
rPAD/7861 PAD:4057 PAD:9765 1.5
rPAD/7862 PAD:4056 PAD:4059 0.0375882
rPAD/7863 PAD:4056 PAD:4057 1.5
rPAD/7864 PAD:4054 PAD:4057 0.0751765
rPAD/7865 PAD:4054 PAD:9762 1.5
rPAD/7866 PAD:4053 PAD:4056 0.0751765
rPAD/7867 PAD:4053 PAD:4054 1.5
rPAD/7868 PAD:4051 PAD:4054 0.0375882
rPAD/7869 PAD:4051 PAD:9759 1.5
rPAD/7870 PAD:4050 PAD:4053 0.0375882
rPAD/7871 PAD:4050 PAD:4051 1.5
rPAD/7872 PAD:4048 PAD:4051 0.0751765
rPAD/7873 PAD:4048 PAD:9756 1.5
rPAD/7874 PAD:4047 PAD:4050 0.0751765
rPAD/7875 PAD:4047 PAD:4048 1.5
rPAD/7876 PAD:4045 PAD:9749 0.0751765
rPAD/7877 PAD:4045 PAD:4048 0.0375882
rPAD/7878 PAD:4045 PAD:9753 1.5
rPAD/7879 PAD:4044 PAD:4047 0.0375882
rPAD/7880 PAD:4044 PAD:4045 1.5
rPAD/7881 PAD:4041 PAD:4044 0.0751765
rPAD/7882 PAD:4041 PAD:9749 1.5
rPAD/7883 PAD:4039 PAD:9749 0.0375882
rPAD/7884 PAD:4039 PAD:9747 1.5
rPAD/7885 PAD:4038 PAD:4041 0.0375882
rPAD/7886 PAD:4038 PAD:4039 1.5
rPAD/7887 PAD:4036 PAD:4039 0.0751765
rPAD/7888 PAD:4036 PAD:9744 1.5
rPAD/7889 PAD:4035 PAD:4038 0.0751765
rPAD/7890 PAD:4035 PAD:4036 1.5
rPAD/7891 PAD:4033 PAD:9737 0.0751765
rPAD/7892 PAD:4033 PAD:4036 0.0375882
rPAD/7893 PAD:4033 PAD:9741 1.5
rPAD/7894 PAD:4032 PAD:4035 0.0375882
rPAD/7895 PAD:4032 PAD:4033 1.5
rPAD/7896 PAD:4029 PAD:4032 0.0751765
rPAD/7897 PAD:4029 PAD:9737 1.5
rPAD/7898 PAD:4026 PAD:4029 0.0375882
rPAD/7899 PAD:4026 PAD:9734 1.5
rPAD/7900 PAD:4023 PAD:4026 0.0751765
rPAD/7901 PAD:4023 PAD:9731 1.5
rPAD/7902 PAD:4020 PAD:4023 0.0375882
rPAD/7903 PAD:4020 PAD:9728 1.5
rPAD/7904 PAD:4017 PAD:4020 0.0751765
rPAD/7905 PAD:4017 PAD:9725 1.5
rPAD/7906 PAD:4015 PAD:9725 0.0375882
rPAD/7907 PAD:4015 PAD:9723 1.5
rPAD/7908 PAD:4014 PAD:4017 0.0375882
rPAD/7909 PAD:4014 PAD:4015 1.5
rPAD/7910 PAD:4012 PAD:9716 0.0375882
rPAD/7911 PAD:4012 PAD:4015 0.0751765
rPAD/7912 PAD:4012 PAD:9720 1.5
rPAD/7913 PAD:4011 PAD:4014 0.0751765
rPAD/7914 PAD:4011 PAD:4012 1.5
rPAD/7915 PAD:4008 PAD:4011 0.0375882
rPAD/7916 PAD:4008 PAD:9716 1.5
rPAD/7917 PAD:4006 PAD:9716 0.0751765
rPAD/7918 PAD:4006 PAD:9714 1.5
rPAD/7919 PAD:4005 PAD:4008 0.0751765
rPAD/7920 PAD:4005 PAD:4006 1.5
rPAD/7921 PAD:4003 PAD:4006 0.0375882
rPAD/7922 PAD:4003 PAD:9711 1.5
rPAD/7923 PAD:4002 PAD:4005 0.0375882
rPAD/7924 PAD:4002 PAD:4003 1.5
rPAD/7925 PAD:4000 PAD:4003 0.0751765
rPAD/7926 PAD:4000 PAD:9708 1.5
rPAD/7927 PAD:3999 PAD:4002 0.0751765
rPAD/7928 PAD:3999 PAD:4000 1.5
rPAD/7929 PAD:3997 PAD:4000 0.0375882
rPAD/7930 PAD:3997 PAD:9705 1.5
rPAD/7931 PAD:3996 PAD:3999 0.0375882
rPAD/7932 PAD:3996 PAD:3997 1.5
rPAD/7933 PAD:3994 PAD:3997 0.0751765
rPAD/7934 PAD:3994 PAD:9702 1.5
rPAD/7935 PAD:3993 PAD:3996 0.0751765
rPAD/7936 PAD:3993 PAD:3994 1.5
rPAD/7937 PAD:3991 PAD:9695 0.0751765
rPAD/7938 PAD:3991 PAD:3994 0.0375882
rPAD/7939 PAD:3991 PAD:9699 1.5
rPAD/7940 PAD:3990 PAD:3993 0.0375882
rPAD/7941 PAD:3990 PAD:3991 1.5
rPAD/7942 PAD:3987 PAD:3990 0.0751765
rPAD/7943 PAD:3987 PAD:9695 1.5
rPAD/7944 PAD:3985 PAD:9695 0.0375882
rPAD/7945 PAD:3985 PAD:9693 1.5
rPAD/7946 PAD:3984 PAD:3987 0.0375882
rPAD/7947 PAD:3984 PAD:3985 1.5
rPAD/7948 PAD:3982 PAD:3985 0.0751765
rPAD/7949 PAD:3982 PAD:9690 1.5
rPAD/7950 PAD:3981 PAD:3984 0.0751765
rPAD/7951 PAD:3981 PAD:3982 1.5
rPAD/7952 PAD:3979 PAD:3982 0.0375882
rPAD/7953 PAD:3979 PAD:9687 1.5
rPAD/7954 PAD:3978 PAD:3981 0.0375882
rPAD/7955 PAD:3978 PAD:3979 1.5
rPAD/7956 PAD:3976 PAD:3979 0.0751765
rPAD/7957 PAD:3976 PAD:9684 1.5
rPAD/7958 PAD:3975 PAD:3978 0.0751765
rPAD/7959 PAD:3975 PAD:3976 1.5
rPAD/7960 PAD:3973 PAD:3976 0.0375882
rPAD/7961 PAD:3973 PAD:9681 1.5
rPAD/7962 PAD:3972 PAD:3975 0.0375882
rPAD/7963 PAD:3972 PAD:3973 1.5
rPAD/7964 PAD:3970 PAD:3973 0.0751765
rPAD/7965 PAD:3970 PAD:9678 1.5
rPAD/7966 PAD:3969 PAD:3972 0.0751765
rPAD/7967 PAD:3969 PAD:3970 1.5
rPAD/7968 PAD:3967 PAD:3970 0.0375882
rPAD/7969 PAD:3967 PAD:9675 1.5
rPAD/7970 PAD:3966 PAD:3969 0.0375882
rPAD/7971 PAD:3966 PAD:3967 1.5
rPAD/7972 PAD:3964 PAD:14833 0.0283817
rPAD/7973 PAD:3964 PAD:3967 0.0751765
rPAD/7974 PAD:3964 PAD:9672 1.5
rPAD/7975 PAD:3963 PAD:9104 0.0378785
rPAD/7976 PAD:3963 PAD:3966 0.0751765
rPAD/7977 PAD:3963 PAD:3964 1.5
rPAD/7978 PAD:3959 PAD:9451 0.0137718
rPAD/7979 PAD:3959 PAD:15014 0.0188456
rPAD/7980 PAD:3958 PAD:3959 2.25
rPAD/7981 PAD:3956 PAD:9451 0.012825
rPAD/7982 PAD:3955 PAD:3958 0.01395
rPAD/7983 PAD:3955 PAD:3956 0.586956
rPAD/7984 PAD:3953 PAD:3956 0.01395
rPAD/7985 PAD:3953 PAD:9666 0.225
rPAD/7986 PAD:3952 PAD:3955 0.01395
rPAD/7987 PAD:3952 PAD:3953 0.586956
rPAD/7988 PAD:3950 PAD:3953 0.0279
rPAD/7989 PAD:3950 PAD:9663 0.586956
rPAD/7990 PAD:3949 PAD:3952 0.0279
rPAD/7991 PAD:3949 PAD:3950 0.586956
rPAD/7992 PAD:3947 PAD:9658 0.01395
rPAD/7993 PAD:3947 PAD:3950 0.01395
rPAD/7994 PAD:3946 PAD:3949 0.01395
rPAD/7995 PAD:3946 PAD:3947 0.586956
rPAD/7996 PAD:3943 PAD:3946 0.0279
rPAD/7997 PAD:3943 PAD:9655 0.586956
rPAD/7998 PAD:3941 PAD:9651 0.01395
rPAD/7999 PAD:3941 PAD:9655 0.01395
rPAD/8000 PAD:3940 PAD:3943 0.01395
rPAD/8001 PAD:3940 PAD:3941 0.586956
rPAD/8002 PAD:3938 PAD:9647 0.01395
rPAD/8003 PAD:3938 PAD:9651 0.01395
rPAD/8004 PAD:3937 PAD:3940 0.0279
rPAD/8005 PAD:3937 PAD:3938 0.586956
rPAD/8006 PAD:3934 PAD:3937 0.0279
rPAD/8007 PAD:3934 PAD:9644 0.586956
rPAD/8008 PAD:3932 PAD:9640 0.01395
rPAD/8009 PAD:3932 PAD:9644 0.01395
rPAD/8010 PAD:3931 PAD:3934 0.01395
rPAD/8011 PAD:3931 PAD:3932 0.586956
rPAD/8012 PAD:3928 PAD:3931 0.0279
rPAD/8013 PAD:3928 PAD:9637 0.586956
rPAD/8014 PAD:3925 PAD:3928 0.01395
rPAD/8015 PAD:3925 PAD:9634 0.586956
rPAD/8016 PAD:3923 PAD:9630 0.01395
rPAD/8017 PAD:3923 PAD:9634 0.01395
rPAD/8018 PAD:3922 PAD:3925 0.01395
rPAD/8019 PAD:3922 PAD:3923 0.586956
rPAD/8020 PAD:3920 PAD:9626 0.01395
rPAD/8021 PAD:3920 PAD:9630 0.01395
rPAD/8022 PAD:3919 PAD:3922 0.0279
rPAD/8023 PAD:3919 PAD:3920 0.586956
rPAD/8024 PAD:3916 PAD:3919 0.0279
rPAD/8025 PAD:3916 PAD:9623 0.586956
rPAD/8026 PAD:3914 PAD:9619 0.01395
rPAD/8027 PAD:3914 PAD:9623 0.01395
rPAD/8028 PAD:3913 PAD:3916 0.01395
rPAD/8029 PAD:3913 PAD:3914 0.586956
rPAD/8030 PAD:3910 PAD:3913 0.0279
rPAD/8031 PAD:3910 PAD:9616 0.586956
rPAD/8032 PAD:3908 PAD:9612 0.01395
rPAD/8033 PAD:3908 PAD:9616 0.01395
rPAD/8034 PAD:3907 PAD:3910 0.01395
rPAD/8035 PAD:3907 PAD:3908 0.586956
rPAD/8036 PAD:3905 PAD:9612 0.01395
rPAD/8037 PAD:3905 PAD:9610 0.586956
rPAD/8038 PAD:3904 PAD:3907 0.0279
rPAD/8039 PAD:3904 PAD:3905 0.586956
rPAD/8040 PAD:3902 PAD:9605 0.01395
rPAD/8041 PAD:3902 PAD:3905 0.01395
rPAD/8042 PAD:3901 PAD:3904 0.01395
rPAD/8043 PAD:3901 PAD:3902 0.586956
rPAD/8044 PAD:3898 PAD:3901 0.0279
rPAD/8045 PAD:3898 PAD:9602 0.586956
rPAD/8046 PAD:3896 PAD:9598 0.01395
rPAD/8047 PAD:3896 PAD:9602 0.01395
rPAD/8048 PAD:3895 PAD:3898 0.01395
rPAD/8049 PAD:3895 PAD:3896 0.586956
rPAD/8050 PAD:3893 PAD:9594 0.01395
rPAD/8051 PAD:3893 PAD:9598 0.01395
rPAD/8052 PAD:3892 PAD:3895 0.0279
rPAD/8053 PAD:3892 PAD:3893 0.586956
rPAD/8054 PAD:3889 PAD:3892 0.0279
rPAD/8055 PAD:3889 PAD:9591 0.586956
rPAD/8056 PAD:3887 PAD:9587 0.01395
rPAD/8057 PAD:3887 PAD:9591 0.01395
rPAD/8058 PAD:3886 PAD:3889 0.01395
rPAD/8059 PAD:3886 PAD:3887 0.586956
rPAD/8060 PAD:3883 PAD:3886 0.0279
rPAD/8061 PAD:3883 PAD:9584 0.586956
rPAD/8062 PAD:3880 PAD:3883 0.01395
rPAD/8063 PAD:3880 PAD:9581 0.586956
rPAD/8064 PAD:3878 PAD:9577 0.01395
rPAD/8065 PAD:3878 PAD:9581 0.01395
rPAD/8066 PAD:3877 PAD:3880 0.01395
rPAD/8067 PAD:3877 PAD:3878 0.586956
rPAD/8068 PAD:3875 PAD:9573 0.01395
rPAD/8069 PAD:3875 PAD:9577 0.01395
rPAD/8070 PAD:3874 PAD:3877 0.0279
rPAD/8071 PAD:3874 PAD:3875 0.586956
rPAD/8072 PAD:3871 PAD:3874 0.0279
rPAD/8073 PAD:3871 PAD:9570 0.586956
rPAD/8074 PAD:3869 PAD:9566 0.01395
rPAD/8075 PAD:3869 PAD:9570 0.01395
rPAD/8076 PAD:3868 PAD:3871 0.01395
rPAD/8077 PAD:3868 PAD:3869 0.586956
rPAD/8078 PAD:3865 PAD:3868 0.0279
rPAD/8079 PAD:3865 PAD:9563 0.586956
rPAD/8080 PAD:3863 PAD:9559 0.01395
rPAD/8081 PAD:3863 PAD:9563 0.01395
rPAD/8082 PAD:3862 PAD:3865 0.01395
rPAD/8083 PAD:3862 PAD:3863 0.586956
rPAD/8084 PAD:3860 PAD:9559 0.01395
rPAD/8085 PAD:3859 PAD:3862 0.0279
rPAD/8086 PAD:3859 PAD:3860 0.586956
rPAD/8087 PAD:3857 PAD:9552 0.01395
rPAD/8088 PAD:3857 PAD:3860 0.01395
rPAD/8089 PAD:3856 PAD:3859 0.01395
rPAD/8090 PAD:3856 PAD:3857 0.586956
rPAD/8091 PAD:3853 PAD:3856 0.0279
rPAD/8092 PAD:3853 PAD:9549 0.586956
rPAD/8093 PAD:3851 PAD:9545 0.01395
rPAD/8094 PAD:3851 PAD:9549 0.01395
rPAD/8095 PAD:3850 PAD:3853 0.01395
rPAD/8096 PAD:3850 PAD:3851 0.586956
rPAD/8097 PAD:3848 PAD:9541 0.01395
rPAD/8098 PAD:3848 PAD:9545 0.01395
rPAD/8099 PAD:3847 PAD:3850 0.0279
rPAD/8100 PAD:3847 PAD:3848 0.586956
rPAD/8101 PAD:3844 PAD:3847 0.0279
rPAD/8102 PAD:3844 PAD:9538 0.586956
rPAD/8103 PAD:3842 PAD:9534 0.01395
rPAD/8104 PAD:3842 PAD:9538 0.01395
rPAD/8105 PAD:3841 PAD:3844 0.01395
rPAD/8106 PAD:3841 PAD:3842 0.586956
rPAD/8107 PAD:3838 PAD:3841 0.0279
rPAD/8108 PAD:3838 PAD:9531 0.586956
rPAD/8109 PAD:3835 PAD:3838 0.01395
rPAD/8110 PAD:3835 PAD:9528 0.586956
rPAD/8111 PAD:3833 PAD:9524 0.01395
rPAD/8112 PAD:3833 PAD:9528 0.01395
rPAD/8113 PAD:3832 PAD:3835 0.01395
rPAD/8114 PAD:3832 PAD:3833 0.586956
rPAD/8115 PAD:3830 PAD:9520 0.01395
rPAD/8116 PAD:3830 PAD:9524 0.01395
rPAD/8117 PAD:3829 PAD:3832 0.0279
rPAD/8118 PAD:3829 PAD:3830 0.586956
rPAD/8119 PAD:3826 PAD:3829 0.0279
rPAD/8120 PAD:3826 PAD:9517 0.586956
rPAD/8121 PAD:3824 PAD:9513 0.01395
rPAD/8122 PAD:3824 PAD:9517 0.01395
rPAD/8123 PAD:3823 PAD:3826 0.01395
rPAD/8124 PAD:3823 PAD:3824 0.586956
rPAD/8125 PAD:3820 PAD:3823 0.0279
rPAD/8126 PAD:3820 PAD:9510 0.586956
rPAD/8127 PAD:3818 PAD:9506 0.01395
rPAD/8128 PAD:3818 PAD:9510 0.01395
rPAD/8129 PAD:3817 PAD:3820 0.01395
rPAD/8130 PAD:3817 PAD:3818 0.586956
rPAD/8131 PAD:3815 PAD:9506 0.01395
rPAD/8132 PAD:3814 PAD:3817 0.0279
rPAD/8133 PAD:3814 PAD:3815 0.586956
rPAD/8134 PAD:3812 PAD:9499 0.01395
rPAD/8135 PAD:3812 PAD:3815 0.01395
rPAD/8136 PAD:3811 PAD:3814 0.01395
rPAD/8137 PAD:3811 PAD:3812 0.586956
rPAD/8138 PAD:3808 PAD:3811 0.0279
rPAD/8139 PAD:3808 PAD:9496 0.586956
rPAD/8140 PAD:3806 PAD:9492 0.01395
rPAD/8141 PAD:3806 PAD:9496 0.01395
rPAD/8142 PAD:3805 PAD:3808 0.01395
rPAD/8143 PAD:3805 PAD:3806 0.586956
rPAD/8144 PAD:3803 PAD:9488 0.01395
rPAD/8145 PAD:3803 PAD:9492 0.01395
rPAD/8146 PAD:3802 PAD:3805 0.0279
rPAD/8147 PAD:3802 PAD:3803 0.586956
rPAD/8148 PAD:3799 PAD:3802 0.0279
rPAD/8149 PAD:3799 PAD:9485 0.586956
rPAD/8150 PAD:3797 PAD:9481 0.01395
rPAD/8151 PAD:3797 PAD:9485 0.01395
rPAD/8152 PAD:3796 PAD:3799 0.01395
rPAD/8153 PAD:3796 PAD:3797 0.586956
rPAD/8154 PAD:3793 PAD:3796 0.0279
rPAD/8155 PAD:3793 PAD:9478 0.586956
rPAD/8156 PAD:3790 PAD:3793 0.01395
rPAD/8157 PAD:3790 PAD:9475 0.586956
rPAD/8158 PAD:3788 PAD:9471 0.01395
rPAD/8159 PAD:3788 PAD:9475 0.01395
rPAD/8160 PAD:3787 PAD:3790 0.01395
rPAD/8161 PAD:3787 PAD:3788 0.586956
rPAD/8162 PAD:3785 PAD:9467 0.01395
rPAD/8163 PAD:3785 PAD:9471 0.01395
rPAD/8164 PAD:3784 PAD:3787 0.0279
rPAD/8165 PAD:3784 PAD:3785 0.586956
rPAD/8166 PAD:3781 PAD:3784 0.0279
rPAD/8167 PAD:3781 PAD:9464 0.586956
rPAD/8168 PAD:3779 PAD:9460 0.01395
rPAD/8169 PAD:3779 PAD:9464 0.01395
rPAD/8170 PAD:3778 PAD:3781 0.01395
rPAD/8171 PAD:3778 PAD:3779 0.586956
rPAD/8172 PAD:3775 PAD:3778 0.0279
rPAD/8173 PAD:3775 PAD:9457 0.586956
rPAD/8174 PAD:3773 PAD:9453 0.01395
rPAD/8175 PAD:3773 PAD:9457 0.01395
rPAD/8176 PAD:3772 PAD:3775 0.01395
rPAD/8177 PAD:3772 PAD:3773 0.586956
rPAD/8178 PAD:3769 PAD:3772 0.0279
rPAD/8179 PAD:3769 PAD:9086 0.586956
rPAD/8180 PAD:3767 PAD:15008 0.35952
rPAD/8181 PAD:3767 PAD:3958 0.007875
rPAD/8182 PAD:3767 PAD:9314 0.0353815
rPAD/8183 PAD:3766 PAD:9089 0.03015
rPAD/8184 PAD:3766 PAD:9093 0.02565
rPAD/8185 PAD:3766 PAD:3769 0.002925
rPAD/8186 PAD:3762 PAD:14799 0.586956
rPAD/8187 PAD:3760 PAD:14788 0.586956
rPAD/8188 PAD:3760 PAD:14786 0.01395
rPAD/8189 PAD:3760 PAD:14793 0.0279
rPAD/8190 PAD:3756 PAD:14767 0.586956
rPAD/8191 PAD:3756 PAD:14765 0.01395
rPAD/8192 PAD:3748 PAD:14725 0.586956
rPAD/8193 PAD:3748 PAD:14722 0.0279
rPAD/8194 PAD:3746 PAD:14714 0.586956
rPAD/8195 PAD:3746 PAD:14712 0.01395
rPAD/8196 PAD:3744 PAD:8984 0.586956
rPAD/8197 PAD:3736 PAD:14661 0.586956
rPAD/8198 PAD:3736 PAD:14659 0.01395
rPAD/8199 PAD:3734 PAD:14648 0.0279
rPAD/8200 PAD:3734 PAD:8939 0.586956
rPAD/8201 PAD:3732 PAD:14640 0.586956
rPAD/8202 PAD:3730 PAD:14629 0.586956
rPAD/8203 PAD:3730 PAD:14634 0.0279
rPAD/8204 PAD:3726 PAD:14608 0.586956
rPAD/8205 PAD:3726 PAD:14606 0.01395
rPAD/8206 PAD:3726 PAD:14613 0.0279
rPAD/8207 PAD:3725 PAD:14811 0.586956
rPAD/8208 PAD:3725 PAD:3762 0.586956
rPAD/8209 PAD:3725 PAD:3760 0.586956
rPAD/8210 PAD:3725 PAD:14779 0.586956
rPAD/8211 PAD:3725 PAD:3756 0.586956
rPAD/8212 PAD:3725 PAD:14758 0.586956
rPAD/8213 PAD:3725 PAD:14747 0.586956
rPAD/8214 PAD:3725 PAD:14736 0.586956
rPAD/8215 PAD:3725 PAD:3748 0.586956
rPAD/8216 PAD:3725 PAD:3746 0.586956
rPAD/8217 PAD:3725 PAD:3744 0.586956
rPAD/8218 PAD:3725 PAD:14694 0.586956
rPAD/8219 PAD:3725 PAD:14683 0.586956
rPAD/8220 PAD:3725 PAD:14673 0.586956
rPAD/8221 PAD:3725 PAD:3736 0.586956
rPAD/8222 PAD:3725 PAD:3734 0.586956
rPAD/8223 PAD:3725 PAD:3732 0.586956
rPAD/8224 PAD:3725 PAD:3730 0.586956
rPAD/8225 PAD:3725 PAD:14620 0.586956
rPAD/8226 PAD:3725 PAD:3726 0.586956
rPAD/8227 PAD:3722 PAD:3725 2.44929e-05
rPAD/8228 PAD:3722 PAD:15142 1.5
rPAD/8229 PAD:3719 PAD:3722 0.000355147
rPAD/8230 PAD:3719 PAD:15004 0.9
rPAD/8231 PAD:3715 PAD:14806 0.586956
rPAD/8232 PAD:3715 PAD:14811 0.0279
rPAD/8233 PAD:3713 PAD:14795 0.586956
rPAD/8234 PAD:3713 PAD:14793 0.01395
rPAD/8235 PAD:3713 PAD:3762 0.0279
rPAD/8236 PAD:3709 PAD:14774 0.586956
rPAD/8237 PAD:3709 PAD:14779 0.0279
rPAD/8238 PAD:3703 PAD:14742 0.586956
rPAD/8239 PAD:3703 PAD:14747 0.0279
rPAD/8240 PAD:3701 PAD:14732 0.586956
rPAD/8241 PAD:3701 PAD:14736 0.01395
rPAD/8242 PAD:3695 PAD:14700 0.586956
rPAD/8243 PAD:3695 PAD:3744 0.0279
rPAD/8244 PAD:3691 PAD:14679 0.586956
rPAD/8245 PAD:3691 PAD:14683 0.01395
rPAD/8246 PAD:3689 PAD:14668 0.586956
rPAD/8247 PAD:3689 PAD:14673 0.0279
rPAD/8248 PAD:3683 PAD:14636 0.586956
rPAD/8249 PAD:3683 PAD:14634 0.01395
rPAD/8250 PAD:3683 PAD:3732 0.0279
rPAD/8251 PAD:3681 PAD:14626 0.586956
rPAD/8252 PAD:3681 PAD:14624 0.01395
rPAD/8253 PAD:3681 PAD:3730 0.01395
rPAD/8254 PAD:3679 PAD:14615 0.586956
rPAD/8255 PAD:3679 PAD:14613 0.01395
rPAD/8256 PAD:3679 PAD:14620 0.0279
rPAD/8257 PAD:3675 PAD:16889 0.000393013
rPAD/8258 PAD:3675 PAD:15000 0.9
rPAD/8259 PAD:3675 PAD:15004 0.0243668
rPAD/8260 PAD:3674 PAD:3719 0.00037964
rPAD/8261 PAD:3674 PAD:14814 0.225
rPAD/8262 PAD:3674 PAD:3715 0.586956
rPAD/8263 PAD:3674 PAD:3713 0.586956
rPAD/8264 PAD:3674 PAD:14786 0.586956
rPAD/8265 PAD:3674 PAD:3709 0.586956
rPAD/8266 PAD:3674 PAD:14765 0.586956
rPAD/8267 PAD:3674 PAD:14754 0.586956
rPAD/8268 PAD:3674 PAD:3703 0.586956
rPAD/8269 PAD:3674 PAD:3701 0.586956
rPAD/8270 PAD:3674 PAD:14722 0.586956
rPAD/8271 PAD:3674 PAD:14712 0.586956
rPAD/8272 PAD:3674 PAD:3695 0.586956
rPAD/8273 PAD:3674 PAD:14690 0.586956
rPAD/8274 PAD:3674 PAD:3691 0.586956
rPAD/8275 PAD:3674 PAD:3689 0.586956
rPAD/8276 PAD:3674 PAD:14659 0.586956
rPAD/8277 PAD:3674 PAD:14648 0.586956
rPAD/8278 PAD:3674 PAD:3683 0.586956
rPAD/8279 PAD:3674 PAD:3681 0.586956
rPAD/8280 PAD:3674 PAD:3679 0.586956
rPAD/8281 PAD:3674 PAD:14606 0.586956
rPAD/8282 PAD:3674 PAD:3675 0.9
rPAD/8283 PAD:3671 PAD:3674 2.44929e-05
rPAD/8284 PAD:3671 PAD:15137 0.346154
rPAD/8285 PAD:3669 PAD:14803 0.586956
rPAD/8286 PAD:3669 PAD:3762 0.0279
rPAD/8287 PAD:3669 PAD:3715 0.01395
rPAD/8288 PAD:3665 PAD:14782 0.586956
rPAD/8289 PAD:3665 PAD:14779 0.0279
rPAD/8290 PAD:3665 PAD:14786 0.01395
rPAD/8291 PAD:3663 PAD:14771 0.586956
rPAD/8292 PAD:3663 PAD:3756 0.0279
rPAD/8293 PAD:3663 PAD:3709 0.01395
rPAD/8294 PAD:3657 PAD:14739 0.586956
rPAD/8295 PAD:3657 PAD:14736 0.0279
rPAD/8296 PAD:3657 PAD:3703 0.01395
rPAD/8297 PAD:3655 PAD:14729 0.586956
rPAD/8298 PAD:3655 PAD:3748 0.0279
rPAD/8299 PAD:3655 PAD:3701 0.01395
rPAD/8300 PAD:3653 PAD:14718 0.586956
rPAD/8301 PAD:3653 PAD:3746 0.0279
rPAD/8302 PAD:3653 PAD:14722 0.01395
rPAD/8303 PAD:3651 PAD:14707 0.586956
rPAD/8304 PAD:3651 PAD:3744 0.01395
rPAD/8305 PAD:3651 PAD:14712 0.0279
rPAD/8306 PAD:3649 PAD:14697 0.586956
rPAD/8307 PAD:3649 PAD:14694 0.0279
rPAD/8308 PAD:3649 PAD:3695 0.01395
rPAD/8309 PAD:3647 PAD:14686 0.586956
rPAD/8310 PAD:3647 PAD:14683 0.0279
rPAD/8311 PAD:3647 PAD:14690 0.01395
rPAD/8312 PAD:3645 PAD:14676 0.586956
rPAD/8313 PAD:3645 PAD:14673 0.0279
rPAD/8314 PAD:3645 PAD:3691 0.01395
rPAD/8315 PAD:3643 PAD:14665 0.586956
rPAD/8316 PAD:3643 PAD:3736 0.0279
rPAD/8317 PAD:3643 PAD:3689 0.01395
rPAD/8318 PAD:3641 PAD:14654 0.586956
rPAD/8319 PAD:3641 PAD:3734 0.01395
rPAD/8320 PAD:3641 PAD:14659 0.0279
rPAD/8321 PAD:3639 PAD:14644 0.586956
rPAD/8322 PAD:3639 PAD:3732 0.0279
rPAD/8323 PAD:3639 PAD:14648 0.01395
rPAD/8324 PAD:3629 PAD:9297 0.9
rPAD/8325 PAD:3629 PAD:16889 0.0483406
rPAD/8326 PAD:3628 PAD:3671 0.000734788
rPAD/8327 PAD:3628 PAD:3669 0.586956
rPAD/8328 PAD:3628 PAD:14793 0.586956
rPAD/8329 PAD:3628 PAD:3665 0.586956
rPAD/8330 PAD:3628 PAD:3663 0.586956
rPAD/8331 PAD:3628 PAD:14761 0.586956
rPAD/8332 PAD:3628 PAD:14751 0.586956
rPAD/8333 PAD:3628 PAD:3657 0.586956
rPAD/8334 PAD:3628 PAD:3655 0.586956
rPAD/8335 PAD:3628 PAD:3653 0.586956
rPAD/8336 PAD:3628 PAD:3651 0.586956
rPAD/8337 PAD:3628 PAD:3649 0.586956
rPAD/8338 PAD:3628 PAD:3647 0.586956
rPAD/8339 PAD:3628 PAD:3645 0.586956
rPAD/8340 PAD:3628 PAD:3643 0.586956
rPAD/8341 PAD:3628 PAD:3641 0.586956
rPAD/8342 PAD:3628 PAD:3639 0.586956
rPAD/8343 PAD:3628 PAD:14634 0.586956
rPAD/8344 PAD:3628 PAD:14624 0.586956
rPAD/8345 PAD:3628 PAD:14613 0.586956
rPAD/8346 PAD:3628 PAD:14602 0.586956
rPAD/8347 PAD:3628 PAD:3629 0.9
rPAD/8348 PAD:3625 PAD:3628 0.000783773
rPAD/8349 PAD:3625 PAD:15134 0.346154
rPAD/8350 PAD:3623 PAD:17018 0.0375328
rPAD/8351 PAD:3623 PAD:14992 0.9
rPAD/8352 PAD:3623 PAD:3629 0.0638646
rPAD/8353 PAD:3622 PAD:3625 0.000211251
rPAD/8354 PAD:3622 PAD:3623 0.9
rPAD/8355 PAD:3614 PAD:14587 1.5
rPAD/8356 PAD:3614 PAD:14585 0.0375882
rPAD/8357 PAD:3614 PAD:14591 0.0751765
rPAD/8358 PAD:3590 PAD:14551 1.5
rPAD/8359 PAD:3590 PAD:14549 0.0375882
rPAD/8360 PAD:3590 PAD:14555 0.0751765
rPAD/8361 PAD:3586 PAD:14545 1.5
rPAD/8362 PAD:3586 PAD:14549 0.0751765
rPAD/8363 PAD:3584 PAD:14542 1.5
rPAD/8364 PAD:3584 PAD:3586 0.0375882
rPAD/8365 PAD:3582 PAD:14539 1.5
rPAD/8366 PAD:3582 PAD:14537 0.0375882
rPAD/8367 PAD:3582 PAD:3584 0.0751765
rPAD/8368 PAD:3578 PAD:14533 1.5
rPAD/8369 PAD:3578 PAD:14537 0.0751765
rPAD/8370 PAD:3576 PAD:14530 1.5
rPAD/8371 PAD:3576 PAD:14528 0.0751765
rPAD/8372 PAD:3576 PAD:3578 0.0375882
rPAD/8373 PAD:3562 PAD:14509 1.5
rPAD/8374 PAD:3562 PAD:14507 0.0375882
rPAD/8375 PAD:3562 PAD:14513 0.0751765
rPAD/8376 PAD:3554 PAD:14497 1.5
rPAD/8377 PAD:3554 PAD:14501 0.0751765
rPAD/8378 PAD:3552 PAD:14494 1.5
rPAD/8379 PAD:3552 PAD:3554 0.0375882
rPAD/8380 PAD:3550 PAD:14491 1.5
rPAD/8381 PAD:3550 PAD:3552 0.0751765
rPAD/8382 PAD:3548 PAD:14488 1.5
rPAD/8383 PAD:3548 PAD:3550 0.0375882
rPAD/8384 PAD:3546 PAD:14485 1.5
rPAD/8385 PAD:3546 PAD:14483 0.0375882
rPAD/8386 PAD:3546 PAD:3548 0.0751765
rPAD/8387 PAD:3540 PAD:14476 1.5
rPAD/8388 PAD:3540 PAD:14474 0.0751765
rPAD/8389 PAD:3540 PAD:14480 0.0375882
rPAD/8390 PAD:3526 PAD:14455 1.5
rPAD/8391 PAD:3526 PAD:14453 0.0375882
rPAD/8392 PAD:3526 PAD:14459 0.0751765
rPAD/8393 PAD:3509 PAD:3622 0.00079602
rPAD/8394 PAD:3509 PAD:14597 1.5
rPAD/8395 PAD:3509 PAD:14594 1.5
rPAD/8396 PAD:3509 PAD:14591 1.5
rPAD/8397 PAD:3509 PAD:3614 1.5
rPAD/8398 PAD:3509 PAD:14585 1.5
rPAD/8399 PAD:3509 PAD:14582 1.5
rPAD/8400 PAD:3509 PAD:14579 1.5
rPAD/8401 PAD:3509 PAD:14576 1.5
rPAD/8402 PAD:3509 PAD:14573 1.5
rPAD/8403 PAD:3509 PAD:14570 1.5
rPAD/8404 PAD:3509 PAD:14567 1.5
rPAD/8405 PAD:3509 PAD:14564 1.5
rPAD/8406 PAD:3509 PAD:14561 1.5
rPAD/8407 PAD:3509 PAD:14558 1.5
rPAD/8408 PAD:3509 PAD:14555 1.5
rPAD/8409 PAD:3509 PAD:3590 1.5
rPAD/8410 PAD:3509 PAD:14549 1.5
rPAD/8411 PAD:3509 PAD:3586 1.5
rPAD/8412 PAD:3509 PAD:3584 1.5
rPAD/8413 PAD:3509 PAD:3582 1.5
rPAD/8414 PAD:3509 PAD:14537 1.5
rPAD/8415 PAD:3509 PAD:3578 1.5
rPAD/8416 PAD:3509 PAD:3576 1.5
rPAD/8417 PAD:3509 PAD:14528 1.5
rPAD/8418 PAD:3509 PAD:14525 1.5
rPAD/8419 PAD:3509 PAD:14522 1.5
rPAD/8420 PAD:3509 PAD:14519 1.5
rPAD/8421 PAD:3509 PAD:14516 1.5
rPAD/8422 PAD:3509 PAD:14513 1.5
rPAD/8423 PAD:3509 PAD:3562 1.5
rPAD/8424 PAD:3509 PAD:14507 1.5
rPAD/8425 PAD:3509 PAD:14504 1.5
rPAD/8426 PAD:3509 PAD:14501 1.5
rPAD/8427 PAD:3509 PAD:3554 1.5
rPAD/8428 PAD:3509 PAD:3552 1.5
rPAD/8429 PAD:3509 PAD:3550 1.5
rPAD/8430 PAD:3509 PAD:3548 1.5
rPAD/8431 PAD:3509 PAD:3546 1.5
rPAD/8432 PAD:3509 PAD:14483 1.5
rPAD/8433 PAD:3509 PAD:14480 1.5
rPAD/8434 PAD:3509 PAD:3540 1.5
rPAD/8435 PAD:3509 PAD:14474 1.5
rPAD/8436 PAD:3509 PAD:14471 1.5
rPAD/8437 PAD:3509 PAD:14468 1.5
rPAD/8438 PAD:3509 PAD:14465 1.5
rPAD/8439 PAD:3509 PAD:14462 1.5
rPAD/8440 PAD:3509 PAD:14459 1.5
rPAD/8441 PAD:3509 PAD:3526 1.5
rPAD/8442 PAD:3509 PAD:14453 1.5
rPAD/8443 PAD:3509 PAD:14450 1.5
rPAD/8444 PAD:3509 PAD:14447 1.5
rPAD/8445 PAD:3509 PAD:14444 1.5
rPAD/8446 PAD:3509 PAD:14441 1.5
rPAD/8447 PAD:3509 PAD:14438 1.5
rPAD/8448 PAD:3509 PAD:14435 1.5
rPAD/8449 PAD:3509 PAD:14432 1.5
rPAD/8450 PAD:3507 PAD:17016 0.0603275
rPAD/8451 PAD:3507 PAD:14987 0.9
rPAD/8452 PAD:3507 PAD:17018 0.0182751
rPAD/8453 PAD:3506 PAD:3509 7.34788e-05
rPAD/8454 PAD:3506 PAD:3507 0.9
rPAD/8455 PAD:3503 PAD:3506 5.81707e-05
rPAD/8456 PAD:3503 PAD:15130 0.346154
rPAD/8457 PAD:3495 PAD:14417 1.5
rPAD/8458 PAD:3495 PAD:14415 0.0375882
rPAD/8459 PAD:3495 PAD:14421 0.0751765
rPAD/8460 PAD:3471 PAD:14381 1.5
rPAD/8461 PAD:3471 PAD:14379 0.0375882
rPAD/8462 PAD:3471 PAD:14385 0.0751765
rPAD/8463 PAD:3467 PAD:14375 1.5
rPAD/8464 PAD:3467 PAD:14379 0.0751765
rPAD/8465 PAD:3465 PAD:14372 1.5
rPAD/8466 PAD:3465 PAD:3467 0.0375882
rPAD/8467 PAD:3463 PAD:14369 1.5
rPAD/8468 PAD:3463 PAD:14367 0.0375882
rPAD/8469 PAD:3463 PAD:3465 0.0751765
rPAD/8470 PAD:3459 PAD:14363 1.5
rPAD/8471 PAD:3459 PAD:14367 0.0751765
rPAD/8472 PAD:3457 PAD:14360 1.5
rPAD/8473 PAD:3457 PAD:14358 0.0751765
rPAD/8474 PAD:3457 PAD:3459 0.0375882
rPAD/8475 PAD:3443 PAD:14339 1.5
rPAD/8476 PAD:3443 PAD:14337 0.0375882
rPAD/8477 PAD:3443 PAD:14343 0.0751765
rPAD/8478 PAD:3435 PAD:14327 1.5
rPAD/8479 PAD:3435 PAD:14331 0.0751765
rPAD/8480 PAD:3433 PAD:14324 1.5
rPAD/8481 PAD:3433 PAD:3435 0.0375882
rPAD/8482 PAD:3431 PAD:14321 1.5
rPAD/8483 PAD:3431 PAD:3433 0.0751765
rPAD/8484 PAD:3429 PAD:14318 1.5
rPAD/8485 PAD:3429 PAD:3431 0.0375882
rPAD/8486 PAD:3427 PAD:14315 1.5
rPAD/8487 PAD:3427 PAD:14313 0.0375882
rPAD/8488 PAD:3427 PAD:3429 0.0751765
rPAD/8489 PAD:3421 PAD:14306 1.5
rPAD/8490 PAD:3421 PAD:14304 0.0751765
rPAD/8491 PAD:3421 PAD:14310 0.0375882
rPAD/8492 PAD:3407 PAD:14285 1.5
rPAD/8493 PAD:3407 PAD:14283 0.0375882
rPAD/8494 PAD:3407 PAD:14289 0.0751765
rPAD/8495 PAD:3390 PAD:3503 0.0011083
rPAD/8496 PAD:3390 PAD:14427 1.5
rPAD/8497 PAD:3390 PAD:14424 1.5
rPAD/8498 PAD:3390 PAD:14421 1.5
rPAD/8499 PAD:3390 PAD:3495 1.5
rPAD/8500 PAD:3390 PAD:14415 1.5
rPAD/8501 PAD:3390 PAD:14412 1.5
rPAD/8502 PAD:3390 PAD:14409 1.5
rPAD/8503 PAD:3390 PAD:14406 1.5
rPAD/8504 PAD:3390 PAD:14403 1.5
rPAD/8505 PAD:3390 PAD:14400 1.5
rPAD/8506 PAD:3390 PAD:14397 1.5
rPAD/8507 PAD:3390 PAD:14394 1.5
rPAD/8508 PAD:3390 PAD:14391 1.5
rPAD/8509 PAD:3390 PAD:14388 1.5
rPAD/8510 PAD:3390 PAD:14385 1.5
rPAD/8511 PAD:3390 PAD:3471 1.5
rPAD/8512 PAD:3390 PAD:14379 1.5
rPAD/8513 PAD:3390 PAD:3467 1.5
rPAD/8514 PAD:3390 PAD:3465 1.5
rPAD/8515 PAD:3390 PAD:3463 1.5
rPAD/8516 PAD:3390 PAD:14367 1.5
rPAD/8517 PAD:3390 PAD:3459 1.5
rPAD/8518 PAD:3390 PAD:3457 1.5
rPAD/8519 PAD:3390 PAD:14358 1.5
rPAD/8520 PAD:3390 PAD:14355 1.5
rPAD/8521 PAD:3390 PAD:14352 1.5
rPAD/8522 PAD:3390 PAD:14349 1.5
rPAD/8523 PAD:3390 PAD:14346 1.5
rPAD/8524 PAD:3390 PAD:14343 1.5
rPAD/8525 PAD:3390 PAD:3443 1.5
rPAD/8526 PAD:3390 PAD:14337 1.5
rPAD/8527 PAD:3390 PAD:14334 1.5
rPAD/8528 PAD:3390 PAD:14331 1.5
rPAD/8529 PAD:3390 PAD:3435 1.5
rPAD/8530 PAD:3390 PAD:3433 1.5
rPAD/8531 PAD:3390 PAD:3431 1.5
rPAD/8532 PAD:3390 PAD:3429 1.5
rPAD/8533 PAD:3390 PAD:3427 1.5
rPAD/8534 PAD:3390 PAD:14313 1.5
rPAD/8535 PAD:3390 PAD:14310 1.5
rPAD/8536 PAD:3390 PAD:3421 1.5
rPAD/8537 PAD:3390 PAD:14304 1.5
rPAD/8538 PAD:3390 PAD:14301 1.5
rPAD/8539 PAD:3390 PAD:14298 1.5
rPAD/8540 PAD:3390 PAD:14295 1.5
rPAD/8541 PAD:3390 PAD:14292 1.5
rPAD/8542 PAD:3390 PAD:14289 1.5
rPAD/8543 PAD:3390 PAD:3407 1.5
rPAD/8544 PAD:3390 PAD:14283 1.5
rPAD/8545 PAD:3390 PAD:14280 1.5
rPAD/8546 PAD:3390 PAD:14277 1.5
rPAD/8547 PAD:3390 PAD:14274 1.5
rPAD/8548 PAD:3390 PAD:14271 1.5
rPAD/8549 PAD:3390 PAD:14268 1.5
rPAD/8550 PAD:3390 PAD:14265 1.5
rPAD/8551 PAD:3390 PAD:14262 1.5
rPAD/8552 PAD:3387 PAD:3390 3.06161e-05
rPAD/8553 PAD:3387 PAD:15126 0.346154
rPAD/8554 PAD:3385 PAD:17014 0.0552183
rPAD/8555 PAD:3385 PAD:14981 0.9
rPAD/8556 PAD:3385 PAD:17016 0.0233843
rPAD/8557 PAD:3384 PAD:3387 0.000107157
rPAD/8558 PAD:3384 PAD:3385 0.9
rPAD/8559 PAD:3382 PAD:17012 0.0780131
rPAD/8560 PAD:3382 PAD:9276 0.9
rPAD/8561 PAD:3382 PAD:17014 0.00058952
rPAD/8562 PAD:3381 PAD:3384 0.000869499
rPAD/8563 PAD:3381 PAD:3382 0.9
rPAD/8564 PAD:3379 PAD:16658 0.041557
rPAD/8565 PAD:3379 PAD:15121 0.346154
rPAD/8566 PAD:3379 PAD:16716 0.0067651
rPAD/8567 PAD:3378 PAD:3381 0.000162266
rPAD/8568 PAD:3378 PAD:3379 0.346154
rPAD/8569 PAD:3370 PAD:14247 1.5
rPAD/8570 PAD:3370 PAD:14245 0.0375882
rPAD/8571 PAD:3370 PAD:14251 0.0751765
rPAD/8572 PAD:3346 PAD:14211 1.5
rPAD/8573 PAD:3346 PAD:14209 0.0375882
rPAD/8574 PAD:3346 PAD:14215 0.0751765
rPAD/8575 PAD:3342 PAD:14205 1.5
rPAD/8576 PAD:3342 PAD:14209 0.0751765
rPAD/8577 PAD:3340 PAD:14202 1.5
rPAD/8578 PAD:3340 PAD:3342 0.0375882
rPAD/8579 PAD:3338 PAD:14199 1.5
rPAD/8580 PAD:3338 PAD:14197 0.0375882
rPAD/8581 PAD:3338 PAD:3340 0.0751765
rPAD/8582 PAD:3334 PAD:14193 1.5
rPAD/8583 PAD:3334 PAD:14197 0.0751765
rPAD/8584 PAD:3332 PAD:14190 1.5
rPAD/8585 PAD:3332 PAD:14188 0.0751765
rPAD/8586 PAD:3332 PAD:3334 0.0375882
rPAD/8587 PAD:3318 PAD:14169 1.5
rPAD/8588 PAD:3318 PAD:14167 0.0375882
rPAD/8589 PAD:3318 PAD:14173 0.0751765
rPAD/8590 PAD:3310 PAD:14157 1.5
rPAD/8591 PAD:3310 PAD:14161 0.0751765
rPAD/8592 PAD:3308 PAD:14154 1.5
rPAD/8593 PAD:3308 PAD:3310 0.0375882
rPAD/8594 PAD:3306 PAD:14151 1.5
rPAD/8595 PAD:3306 PAD:3308 0.0751765
rPAD/8596 PAD:3304 PAD:14148 1.5
rPAD/8597 PAD:3304 PAD:3306 0.0375882
rPAD/8598 PAD:3302 PAD:14145 1.5
rPAD/8599 PAD:3302 PAD:14143 0.0375882
rPAD/8600 PAD:3302 PAD:3304 0.0751765
rPAD/8601 PAD:3296 PAD:14136 1.5
rPAD/8602 PAD:3296 PAD:14134 0.0751765
rPAD/8603 PAD:3296 PAD:14140 0.0375882
rPAD/8604 PAD:3282 PAD:14115 1.5
rPAD/8605 PAD:3282 PAD:14113 0.0375882
rPAD/8606 PAD:3282 PAD:14119 0.0751765
rPAD/8607 PAD:3265 PAD:3378 5.51091e-05
rPAD/8608 PAD:3265 PAD:14257 1.5
rPAD/8609 PAD:3265 PAD:14254 1.5
rPAD/8610 PAD:3265 PAD:14251 1.5
rPAD/8611 PAD:3265 PAD:3370 1.5
rPAD/8612 PAD:3265 PAD:14245 1.5
rPAD/8613 PAD:3265 PAD:14242 1.5
rPAD/8614 PAD:3265 PAD:14239 1.5
rPAD/8615 PAD:3265 PAD:14236 1.5
rPAD/8616 PAD:3265 PAD:14233 1.5
rPAD/8617 PAD:3265 PAD:14230 1.5
rPAD/8618 PAD:3265 PAD:14227 1.5
rPAD/8619 PAD:3265 PAD:14224 1.5
rPAD/8620 PAD:3265 PAD:14221 1.5
rPAD/8621 PAD:3265 PAD:14218 1.5
rPAD/8622 PAD:3265 PAD:14215 1.5
rPAD/8623 PAD:3265 PAD:3346 1.5
rPAD/8624 PAD:3265 PAD:14209 1.5
rPAD/8625 PAD:3265 PAD:3342 1.5
rPAD/8626 PAD:3265 PAD:3340 1.5
rPAD/8627 PAD:3265 PAD:3338 1.5
rPAD/8628 PAD:3265 PAD:14197 1.5
rPAD/8629 PAD:3265 PAD:3334 1.5
rPAD/8630 PAD:3265 PAD:3332 1.5
rPAD/8631 PAD:3265 PAD:14188 1.5
rPAD/8632 PAD:3265 PAD:14185 1.5
rPAD/8633 PAD:3265 PAD:14182 1.5
rPAD/8634 PAD:3265 PAD:14179 1.5
rPAD/8635 PAD:3265 PAD:14176 1.5
rPAD/8636 PAD:3265 PAD:14173 1.5
rPAD/8637 PAD:3265 PAD:3318 1.5
rPAD/8638 PAD:3265 PAD:14167 1.5
rPAD/8639 PAD:3265 PAD:14164 1.5
rPAD/8640 PAD:3265 PAD:14161 1.5
rPAD/8641 PAD:3265 PAD:3310 1.5
rPAD/8642 PAD:3265 PAD:3308 1.5
rPAD/8643 PAD:3265 PAD:3306 1.5
rPAD/8644 PAD:3265 PAD:3304 1.5
rPAD/8645 PAD:3265 PAD:3302 1.5
rPAD/8646 PAD:3265 PAD:14143 1.5
rPAD/8647 PAD:3265 PAD:14140 1.5
rPAD/8648 PAD:3265 PAD:3296 1.5
rPAD/8649 PAD:3265 PAD:14134 1.5
rPAD/8650 PAD:3265 PAD:14131 1.5
rPAD/8651 PAD:3265 PAD:14128 1.5
rPAD/8652 PAD:3265 PAD:14125 1.5
rPAD/8653 PAD:3265 PAD:14122 1.5
rPAD/8654 PAD:3265 PAD:14119 1.5
rPAD/8655 PAD:3265 PAD:3282 1.5
rPAD/8656 PAD:3265 PAD:14113 1.5
rPAD/8657 PAD:3265 PAD:14110 1.5
rPAD/8658 PAD:3265 PAD:14107 1.5
rPAD/8659 PAD:3265 PAD:14104 1.5
rPAD/8660 PAD:3265 PAD:14101 1.5
rPAD/8661 PAD:3265 PAD:14098 1.5
rPAD/8662 PAD:3265 PAD:14095 1.5
rPAD/8663 PAD:3265 PAD:14092 1.5
rPAD/8664 PAD:3263 PAD:14971 0.9
rPAD/8665 PAD:3263 PAD:17012 0.00569869
rPAD/8666 PAD:3262 PAD:3265 0.00108687
rPAD/8667 PAD:3262 PAD:3263 0.9
rPAD/8668 PAD:3254 PAD:14077 1.5
rPAD/8669 PAD:3254 PAD:14075 0.0375882
rPAD/8670 PAD:3254 PAD:14081 0.0751765
rPAD/8671 PAD:3230 PAD:14041 1.5
rPAD/8672 PAD:3230 PAD:14039 0.0375882
rPAD/8673 PAD:3230 PAD:14045 0.0751765
rPAD/8674 PAD:3226 PAD:14035 1.5
rPAD/8675 PAD:3226 PAD:14039 0.0751765
rPAD/8676 PAD:3224 PAD:14032 1.5
rPAD/8677 PAD:3224 PAD:3226 0.0375882
rPAD/8678 PAD:3222 PAD:14029 1.5
rPAD/8679 PAD:3222 PAD:14027 0.0375882
rPAD/8680 PAD:3222 PAD:3224 0.0751765
rPAD/8681 PAD:3218 PAD:14023 1.5
rPAD/8682 PAD:3218 PAD:14027 0.0751765
rPAD/8683 PAD:3216 PAD:14020 1.5
rPAD/8684 PAD:3216 PAD:14018 0.0751765
rPAD/8685 PAD:3216 PAD:3218 0.0375882
rPAD/8686 PAD:3202 PAD:13999 1.5
rPAD/8687 PAD:3202 PAD:13997 0.0375882
rPAD/8688 PAD:3202 PAD:14003 0.0751765
rPAD/8689 PAD:3194 PAD:13987 1.5
rPAD/8690 PAD:3194 PAD:13991 0.0751765
rPAD/8691 PAD:3192 PAD:13984 1.5
rPAD/8692 PAD:3192 PAD:3194 0.0375882
rPAD/8693 PAD:3190 PAD:13981 1.5
rPAD/8694 PAD:3190 PAD:3192 0.0751765
rPAD/8695 PAD:3188 PAD:13978 1.5
rPAD/8696 PAD:3188 PAD:3190 0.0375882
rPAD/8697 PAD:3186 PAD:13975 1.5
rPAD/8698 PAD:3186 PAD:13973 0.0375882
rPAD/8699 PAD:3186 PAD:3188 0.0751765
rPAD/8700 PAD:3180 PAD:13966 1.5
rPAD/8701 PAD:3180 PAD:13964 0.0751765
rPAD/8702 PAD:3180 PAD:13970 0.0375882
rPAD/8703 PAD:3166 PAD:13945 1.5
rPAD/8704 PAD:3166 PAD:13943 0.0375882
rPAD/8705 PAD:3166 PAD:13949 0.0751765
rPAD/8706 PAD:3149 PAD:3262 0.000153081
rPAD/8707 PAD:3149 PAD:14087 1.5
rPAD/8708 PAD:3149 PAD:14084 1.5
rPAD/8709 PAD:3149 PAD:14081 1.5
rPAD/8710 PAD:3149 PAD:3254 1.5
rPAD/8711 PAD:3149 PAD:14075 1.5
rPAD/8712 PAD:3149 PAD:14072 1.5
rPAD/8713 PAD:3149 PAD:14069 1.5
rPAD/8714 PAD:3149 PAD:14066 1.5
rPAD/8715 PAD:3149 PAD:14063 1.5
rPAD/8716 PAD:3149 PAD:14060 1.5
rPAD/8717 PAD:3149 PAD:14057 1.5
rPAD/8718 PAD:3149 PAD:14054 1.5
rPAD/8719 PAD:3149 PAD:14051 1.5
rPAD/8720 PAD:3149 PAD:14048 1.5
rPAD/8721 PAD:3149 PAD:14045 1.5
rPAD/8722 PAD:3149 PAD:3230 1.5
rPAD/8723 PAD:3149 PAD:14039 1.5
rPAD/8724 PAD:3149 PAD:3226 1.5
rPAD/8725 PAD:3149 PAD:3224 1.5
rPAD/8726 PAD:3149 PAD:3222 1.5
rPAD/8727 PAD:3149 PAD:14027 1.5
rPAD/8728 PAD:3149 PAD:3218 1.5
rPAD/8729 PAD:3149 PAD:3216 1.5
rPAD/8730 PAD:3149 PAD:14018 1.5
rPAD/8731 PAD:3149 PAD:14015 1.5
rPAD/8732 PAD:3149 PAD:14012 1.5
rPAD/8733 PAD:3149 PAD:14009 1.5
rPAD/8734 PAD:3149 PAD:14006 1.5
rPAD/8735 PAD:3149 PAD:14003 1.5
rPAD/8736 PAD:3149 PAD:3202 1.5
rPAD/8737 PAD:3149 PAD:13997 1.5
rPAD/8738 PAD:3149 PAD:13994 1.5
rPAD/8739 PAD:3149 PAD:13991 1.5
rPAD/8740 PAD:3149 PAD:3194 1.5
rPAD/8741 PAD:3149 PAD:3192 1.5
rPAD/8742 PAD:3149 PAD:3190 1.5
rPAD/8743 PAD:3149 PAD:3188 1.5
rPAD/8744 PAD:3149 PAD:3186 1.5
rPAD/8745 PAD:3149 PAD:13973 1.5
rPAD/8746 PAD:3149 PAD:13970 1.5
rPAD/8747 PAD:3149 PAD:3180 1.5
rPAD/8748 PAD:3149 PAD:13964 1.5
rPAD/8749 PAD:3149 PAD:13961 1.5
rPAD/8750 PAD:3149 PAD:13958 1.5
rPAD/8751 PAD:3149 PAD:13955 1.5
rPAD/8752 PAD:3149 PAD:13952 1.5
rPAD/8753 PAD:3149 PAD:13949 1.5
rPAD/8754 PAD:3149 PAD:3166 1.5
rPAD/8755 PAD:3149 PAD:13943 1.5
rPAD/8756 PAD:3149 PAD:13940 1.5
rPAD/8757 PAD:3149 PAD:13937 1.5
rPAD/8758 PAD:3149 PAD:13934 1.5
rPAD/8759 PAD:3149 PAD:13931 1.5
rPAD/8760 PAD:3149 PAD:13928 1.5
rPAD/8761 PAD:3149 PAD:13925 1.5
rPAD/8762 PAD:3149 PAD:13922 1.5
rPAD/8763 PAD:3147 PAD:16600 0.0299597
rPAD/8764 PAD:3147 PAD:15117 0.346154
rPAD/8765 PAD:3147 PAD:16658 0.0183624
rPAD/8766 PAD:3146 PAD:3149 0.000223498
rPAD/8767 PAD:3146 PAD:3147 0.346154
rPAD/8768 PAD:3144 PAD:17009 0.0170961
rPAD/8769 PAD:3144 PAD:14968 0.9
rPAD/8770 PAD:3144 PAD:3263 0.0558079
rPAD/8771 PAD:3143 PAD:3146 0.00049292
rPAD/8772 PAD:3143 PAD:3144 0.9
rPAD/8773 PAD:3135 PAD:13907 1.5
rPAD/8774 PAD:3135 PAD:13905 0.0375882
rPAD/8775 PAD:3135 PAD:13911 0.0751765
rPAD/8776 PAD:3111 PAD:13871 1.5
rPAD/8777 PAD:3111 PAD:13869 0.0375882
rPAD/8778 PAD:3111 PAD:13875 0.0751765
rPAD/8779 PAD:3107 PAD:13865 1.5
rPAD/8780 PAD:3107 PAD:13869 0.0751765
rPAD/8781 PAD:3105 PAD:13862 1.5
rPAD/8782 PAD:3105 PAD:3107 0.0375882
rPAD/8783 PAD:3103 PAD:13859 1.5
rPAD/8784 PAD:3103 PAD:13857 0.0375882
rPAD/8785 PAD:3103 PAD:3105 0.0751765
rPAD/8786 PAD:3099 PAD:13853 1.5
rPAD/8787 PAD:3099 PAD:13857 0.0751765
rPAD/8788 PAD:3097 PAD:13850 1.5
rPAD/8789 PAD:3097 PAD:13848 0.0751765
rPAD/8790 PAD:3097 PAD:3099 0.0375882
rPAD/8791 PAD:3083 PAD:13829 1.5
rPAD/8792 PAD:3083 PAD:13827 0.0375882
rPAD/8793 PAD:3083 PAD:13833 0.0751765
rPAD/8794 PAD:3075 PAD:13817 1.5
rPAD/8795 PAD:3075 PAD:13821 0.0751765
rPAD/8796 PAD:3073 PAD:13814 1.5
rPAD/8797 PAD:3073 PAD:3075 0.0375882
rPAD/8798 PAD:3071 PAD:13811 1.5
rPAD/8799 PAD:3071 PAD:3073 0.0751765
rPAD/8800 PAD:3069 PAD:13808 1.5
rPAD/8801 PAD:3069 PAD:3071 0.0375882
rPAD/8802 PAD:3067 PAD:13805 1.5
rPAD/8803 PAD:3067 PAD:13803 0.0375882
rPAD/8804 PAD:3067 PAD:3069 0.0751765
rPAD/8805 PAD:3061 PAD:13796 1.5
rPAD/8806 PAD:3061 PAD:13794 0.0751765
rPAD/8807 PAD:3061 PAD:13800 0.0375882
rPAD/8808 PAD:3047 PAD:13775 1.5
rPAD/8809 PAD:3047 PAD:13773 0.0375882
rPAD/8810 PAD:3047 PAD:13779 0.0751765
rPAD/8811 PAD:3030 PAD:3143 0.000499043
rPAD/8812 PAD:3030 PAD:13917 1.5
rPAD/8813 PAD:3030 PAD:13914 1.5
rPAD/8814 PAD:3030 PAD:13911 1.5
rPAD/8815 PAD:3030 PAD:3135 1.5
rPAD/8816 PAD:3030 PAD:13905 1.5
rPAD/8817 PAD:3030 PAD:13902 1.5
rPAD/8818 PAD:3030 PAD:13899 1.5
rPAD/8819 PAD:3030 PAD:13896 1.5
rPAD/8820 PAD:3030 PAD:13893 1.5
rPAD/8821 PAD:3030 PAD:13890 1.5
rPAD/8822 PAD:3030 PAD:13887 1.5
rPAD/8823 PAD:3030 PAD:13884 1.5
rPAD/8824 PAD:3030 PAD:13881 1.5
rPAD/8825 PAD:3030 PAD:13878 1.5
rPAD/8826 PAD:3030 PAD:13875 1.5
rPAD/8827 PAD:3030 PAD:3111 1.5
rPAD/8828 PAD:3030 PAD:13869 1.5
rPAD/8829 PAD:3030 PAD:3107 1.5
rPAD/8830 PAD:3030 PAD:3105 1.5
rPAD/8831 PAD:3030 PAD:3103 1.5
rPAD/8832 PAD:3030 PAD:13857 1.5
rPAD/8833 PAD:3030 PAD:3099 1.5
rPAD/8834 PAD:3030 PAD:3097 1.5
rPAD/8835 PAD:3030 PAD:13848 1.5
rPAD/8836 PAD:3030 PAD:13845 1.5
rPAD/8837 PAD:3030 PAD:13842 1.5
rPAD/8838 PAD:3030 PAD:13839 1.5
rPAD/8839 PAD:3030 PAD:13836 1.5
rPAD/8840 PAD:3030 PAD:13833 1.5
rPAD/8841 PAD:3030 PAD:3083 1.5
rPAD/8842 PAD:3030 PAD:13827 1.5
rPAD/8843 PAD:3030 PAD:13824 1.5
rPAD/8844 PAD:3030 PAD:13821 1.5
rPAD/8845 PAD:3030 PAD:3075 1.5
rPAD/8846 PAD:3030 PAD:3073 1.5
rPAD/8847 PAD:3030 PAD:3071 1.5
rPAD/8848 PAD:3030 PAD:3069 1.5
rPAD/8849 PAD:3030 PAD:3067 1.5
rPAD/8850 PAD:3030 PAD:13803 1.5
rPAD/8851 PAD:3030 PAD:13800 1.5
rPAD/8852 PAD:3030 PAD:3061 1.5
rPAD/8853 PAD:3030 PAD:13794 1.5
rPAD/8854 PAD:3030 PAD:13791 1.5
rPAD/8855 PAD:3030 PAD:13788 1.5
rPAD/8856 PAD:3030 PAD:13785 1.5
rPAD/8857 PAD:3030 PAD:13782 1.5
rPAD/8858 PAD:3030 PAD:13779 1.5
rPAD/8859 PAD:3030 PAD:3047 1.5
rPAD/8860 PAD:3030 PAD:13773 1.5
rPAD/8861 PAD:3030 PAD:13770 1.5
rPAD/8862 PAD:3030 PAD:13767 1.5
rPAD/8863 PAD:3030 PAD:13764 1.5
rPAD/8864 PAD:3030 PAD:13761 1.5
rPAD/8865 PAD:3030 PAD:13758 1.5
rPAD/8866 PAD:3030 PAD:13755 1.5
rPAD/8867 PAD:3030 PAD:13752 1.5
rPAD/8868 PAD:3028 PAD:16542 0.0333423
rPAD/8869 PAD:3028 PAD:15113 0.346154
rPAD/8870 PAD:3028 PAD:16600 0.0149799
rPAD/8871 PAD:3027 PAD:3030 0.000146958
rPAD/8872 PAD:3027 PAD:3028 0.346154
rPAD/8873 PAD:3025 PAD:17007 0.0119869
rPAD/8874 PAD:3025 PAD:14963 0.9
rPAD/8875 PAD:3025 PAD:17009 0.0666157
rPAD/8876 PAD:3024 PAD:3027 0.000658247
rPAD/8877 PAD:3024 PAD:3025 0.9
rPAD/8878 PAD:3016 PAD:13737 1.5
rPAD/8879 PAD:3016 PAD:13735 0.0375882
rPAD/8880 PAD:3016 PAD:13741 0.0751765
rPAD/8881 PAD:2992 PAD:13701 1.5
rPAD/8882 PAD:2992 PAD:13699 0.0375882
rPAD/8883 PAD:2992 PAD:13705 0.0751765
rPAD/8884 PAD:2988 PAD:13695 1.5
rPAD/8885 PAD:2988 PAD:13699 0.0751765
rPAD/8886 PAD:2986 PAD:13692 1.5
rPAD/8887 PAD:2986 PAD:2988 0.0375882
rPAD/8888 PAD:2984 PAD:13689 1.5
rPAD/8889 PAD:2984 PAD:13687 0.0375882
rPAD/8890 PAD:2984 PAD:2986 0.0751765
rPAD/8891 PAD:2980 PAD:13683 1.5
rPAD/8892 PAD:2980 PAD:13687 0.0751765
rPAD/8893 PAD:2978 PAD:13680 1.5
rPAD/8894 PAD:2978 PAD:13678 0.0751765
rPAD/8895 PAD:2978 PAD:2980 0.0375882
rPAD/8896 PAD:2964 PAD:13659 1.5
rPAD/8897 PAD:2964 PAD:13657 0.0375882
rPAD/8898 PAD:2964 PAD:13663 0.0751765
rPAD/8899 PAD:2956 PAD:13647 1.5
rPAD/8900 PAD:2956 PAD:13651 0.0751765
rPAD/8901 PAD:2954 PAD:13644 1.5
rPAD/8902 PAD:2954 PAD:2956 0.0375882
rPAD/8903 PAD:2952 PAD:13641 1.5
rPAD/8904 PAD:2952 PAD:2954 0.0751765
rPAD/8905 PAD:2950 PAD:13638 1.5
rPAD/8906 PAD:2950 PAD:2952 0.0375882
rPAD/8907 PAD:2948 PAD:13635 1.5
rPAD/8908 PAD:2948 PAD:13633 0.0375882
rPAD/8909 PAD:2948 PAD:2950 0.0751765
rPAD/8910 PAD:2942 PAD:13626 1.5
rPAD/8911 PAD:2942 PAD:13624 0.0751765
rPAD/8912 PAD:2942 PAD:13630 0.0375882
rPAD/8913 PAD:2928 PAD:13605 1.5
rPAD/8914 PAD:2928 PAD:13603 0.0375882
rPAD/8915 PAD:2928 PAD:13609 0.0751765
rPAD/8916 PAD:2911 PAD:3024 0.000419441
rPAD/8917 PAD:2911 PAD:13747 1.5
rPAD/8918 PAD:2911 PAD:13744 1.5
rPAD/8919 PAD:2911 PAD:13741 1.5
rPAD/8920 PAD:2911 PAD:3016 1.5
rPAD/8921 PAD:2911 PAD:13735 1.5
rPAD/8922 PAD:2911 PAD:13732 1.5
rPAD/8923 PAD:2911 PAD:13729 1.5
rPAD/8924 PAD:2911 PAD:13726 1.5
rPAD/8925 PAD:2911 PAD:13723 1.5
rPAD/8926 PAD:2911 PAD:13720 1.5
rPAD/8927 PAD:2911 PAD:13717 1.5
rPAD/8928 PAD:2911 PAD:13714 1.5
rPAD/8929 PAD:2911 PAD:13711 1.5
rPAD/8930 PAD:2911 PAD:13708 1.5
rPAD/8931 PAD:2911 PAD:13705 1.5
rPAD/8932 PAD:2911 PAD:2992 1.5
rPAD/8933 PAD:2911 PAD:13699 1.5
rPAD/8934 PAD:2911 PAD:2988 1.5
rPAD/8935 PAD:2911 PAD:2986 1.5
rPAD/8936 PAD:2911 PAD:2984 1.5
rPAD/8937 PAD:2911 PAD:13687 1.5
rPAD/8938 PAD:2911 PAD:2980 1.5
rPAD/8939 PAD:2911 PAD:2978 1.5
rPAD/8940 PAD:2911 PAD:13678 1.5
rPAD/8941 PAD:2911 PAD:13675 1.5
rPAD/8942 PAD:2911 PAD:13672 1.5
rPAD/8943 PAD:2911 PAD:13669 1.5
rPAD/8944 PAD:2911 PAD:13666 1.5
rPAD/8945 PAD:2911 PAD:13663 1.5
rPAD/8946 PAD:2911 PAD:2964 1.5
rPAD/8947 PAD:2911 PAD:13657 1.5
rPAD/8948 PAD:2911 PAD:13654 1.5
rPAD/8949 PAD:2911 PAD:13651 1.5
rPAD/8950 PAD:2911 PAD:2956 1.5
rPAD/8951 PAD:2911 PAD:2954 1.5
rPAD/8952 PAD:2911 PAD:2952 1.5
rPAD/8953 PAD:2911 PAD:2950 1.5
rPAD/8954 PAD:2911 PAD:2948 1.5
rPAD/8955 PAD:2911 PAD:13633 1.5
rPAD/8956 PAD:2911 PAD:13630 1.5
rPAD/8957 PAD:2911 PAD:2942 1.5
rPAD/8958 PAD:2911 PAD:13624 1.5
rPAD/8959 PAD:2911 PAD:13621 1.5
rPAD/8960 PAD:2911 PAD:13618 1.5
rPAD/8961 PAD:2911 PAD:13615 1.5
rPAD/8962 PAD:2911 PAD:13612 1.5
rPAD/8963 PAD:2911 PAD:13609 1.5
rPAD/8964 PAD:2911 PAD:2928 1.5
rPAD/8965 PAD:2911 PAD:13603 1.5
rPAD/8966 PAD:2911 PAD:13600 1.5
rPAD/8967 PAD:2911 PAD:13597 1.5
rPAD/8968 PAD:2911 PAD:13594 1.5
rPAD/8969 PAD:2911 PAD:13591 1.5
rPAD/8970 PAD:2911 PAD:13588 1.5
rPAD/8971 PAD:2911 PAD:13585 1.5
rPAD/8972 PAD:2911 PAD:13582 1.5
rPAD/8973 PAD:2909 PAD:16484 0.0367248
rPAD/8974 PAD:2909 PAD:15109 0.346154
rPAD/8975 PAD:2909 PAD:16542 0.0115973
rPAD/8976 PAD:2908 PAD:2911 6.12323e-05
rPAD/8977 PAD:2908 PAD:2909 0.346154
rPAD/8978 PAD:2906 PAD:17005 0.0347817
rPAD/8979 PAD:2906 PAD:14958 0.9
rPAD/8980 PAD:2906 PAD:17007 0.043821
rPAD/8981 PAD:2905 PAD:2908 0.000388825
rPAD/8982 PAD:2905 PAD:2906 0.9
rPAD/8983 PAD:2903 PAD:16426 0.0401074
rPAD/8984 PAD:2903 PAD:15105 0.346154
rPAD/8985 PAD:2903 PAD:16484 0.00821477
rPAD/8986 PAD:2902 PAD:2905 0.000750096
rPAD/8987 PAD:2902 PAD:2903 0.346154
rPAD/8988 PAD:2894 PAD:13567 1.5
rPAD/8989 PAD:2894 PAD:13565 0.0375882
rPAD/8990 PAD:2894 PAD:13571 0.0751765
rPAD/8991 PAD:2870 PAD:13531 1.5
rPAD/8992 PAD:2870 PAD:13529 0.0375882
rPAD/8993 PAD:2870 PAD:13535 0.0751765
rPAD/8994 PAD:2866 PAD:13525 1.5
rPAD/8995 PAD:2866 PAD:13529 0.0751765
rPAD/8996 PAD:2864 PAD:13522 1.5
rPAD/8997 PAD:2864 PAD:2866 0.0375882
rPAD/8998 PAD:2862 PAD:13519 1.5
rPAD/8999 PAD:2862 PAD:13517 0.0375882
rPAD/9000 PAD:2862 PAD:2864 0.0751765
rPAD/9001 PAD:2858 PAD:13513 1.5
rPAD/9002 PAD:2858 PAD:13517 0.0751765
rPAD/9003 PAD:2856 PAD:13510 1.5
rPAD/9004 PAD:2856 PAD:13508 0.0751765
rPAD/9005 PAD:2856 PAD:2858 0.0375882
rPAD/9006 PAD:2842 PAD:13489 1.5
rPAD/9007 PAD:2842 PAD:13487 0.0375882
rPAD/9008 PAD:2842 PAD:13493 0.0751765
rPAD/9009 PAD:2834 PAD:13477 1.5
rPAD/9010 PAD:2834 PAD:13481 0.0751765
rPAD/9011 PAD:2832 PAD:13474 1.5
rPAD/9012 PAD:2832 PAD:2834 0.0375882
rPAD/9013 PAD:2830 PAD:13471 1.5
rPAD/9014 PAD:2830 PAD:2832 0.0751765
rPAD/9015 PAD:2828 PAD:13468 1.5
rPAD/9016 PAD:2828 PAD:2830 0.0375882
rPAD/9017 PAD:2826 PAD:13465 1.5
rPAD/9018 PAD:2826 PAD:13463 0.0375882
rPAD/9019 PAD:2826 PAD:2828 0.0751765
rPAD/9020 PAD:2820 PAD:13456 1.5
rPAD/9021 PAD:2820 PAD:13454 0.0751765
rPAD/9022 PAD:2820 PAD:13460 0.0375882
rPAD/9023 PAD:2806 PAD:13435 1.5
rPAD/9024 PAD:2806 PAD:13433 0.0375882
rPAD/9025 PAD:2806 PAD:13439 0.0751765
rPAD/9026 PAD:2789 PAD:2902 1.22465e-05
rPAD/9027 PAD:2789 PAD:13577 1.5
rPAD/9028 PAD:2789 PAD:13574 1.5
rPAD/9029 PAD:2789 PAD:13571 1.5
rPAD/9030 PAD:2789 PAD:2894 1.5
rPAD/9031 PAD:2789 PAD:13565 1.5
rPAD/9032 PAD:2789 PAD:13562 1.5
rPAD/9033 PAD:2789 PAD:13559 1.5
rPAD/9034 PAD:2789 PAD:13556 1.5
rPAD/9035 PAD:2789 PAD:13553 1.5
rPAD/9036 PAD:2789 PAD:13550 1.5
rPAD/9037 PAD:2789 PAD:13547 1.5
rPAD/9038 PAD:2789 PAD:13544 1.5
rPAD/9039 PAD:2789 PAD:13541 1.5
rPAD/9040 PAD:2789 PAD:13538 1.5
rPAD/9041 PAD:2789 PAD:13535 1.5
rPAD/9042 PAD:2789 PAD:2870 1.5
rPAD/9043 PAD:2789 PAD:13529 1.5
rPAD/9044 PAD:2789 PAD:2866 1.5
rPAD/9045 PAD:2789 PAD:2864 1.5
rPAD/9046 PAD:2789 PAD:2862 1.5
rPAD/9047 PAD:2789 PAD:13517 1.5
rPAD/9048 PAD:2789 PAD:2858 1.5
rPAD/9049 PAD:2789 PAD:2856 1.5
rPAD/9050 PAD:2789 PAD:13508 1.5
rPAD/9051 PAD:2789 PAD:13505 1.5
rPAD/9052 PAD:2789 PAD:13502 1.5
rPAD/9053 PAD:2789 PAD:13499 1.5
rPAD/9054 PAD:2789 PAD:13496 1.5
rPAD/9055 PAD:2789 PAD:13493 1.5
rPAD/9056 PAD:2789 PAD:2842 1.5
rPAD/9057 PAD:2789 PAD:13487 1.5
rPAD/9058 PAD:2789 PAD:13484 1.5
rPAD/9059 PAD:2789 PAD:13481 1.5
rPAD/9060 PAD:2789 PAD:2834 1.5
rPAD/9061 PAD:2789 PAD:2832 1.5
rPAD/9062 PAD:2789 PAD:2830 1.5
rPAD/9063 PAD:2789 PAD:2828 1.5
rPAD/9064 PAD:2789 PAD:2826 1.5
rPAD/9065 PAD:2789 PAD:13463 1.5
rPAD/9066 PAD:2789 PAD:13460 1.5
rPAD/9067 PAD:2789 PAD:2820 1.5
rPAD/9068 PAD:2789 PAD:13454 1.5
rPAD/9069 PAD:2789 PAD:13451 1.5
rPAD/9070 PAD:2789 PAD:13448 1.5
rPAD/9071 PAD:2789 PAD:13445 1.5
rPAD/9072 PAD:2789 PAD:13442 1.5
rPAD/9073 PAD:2789 PAD:13439 1.5
rPAD/9074 PAD:2789 PAD:2806 1.5
rPAD/9075 PAD:2789 PAD:13433 1.5
rPAD/9076 PAD:2789 PAD:13430 1.5
rPAD/9077 PAD:2789 PAD:13427 1.5
rPAD/9078 PAD:2789 PAD:13424 1.5
rPAD/9079 PAD:2789 PAD:13421 1.5
rPAD/9080 PAD:2789 PAD:13418 1.5
rPAD/9081 PAD:2789 PAD:13415 1.5
rPAD/9082 PAD:2789 PAD:13412 1.5
rPAD/9083 PAD:2787 PAD:17003 0.0296725
rPAD/9084 PAD:2787 PAD:14952 0.9
rPAD/9085 PAD:2787 PAD:17005 0.0489301
rPAD/9086 PAD:2786 PAD:2789 0.000541906
rPAD/9087 PAD:2786 PAD:2787 0.9
rPAD/9088 PAD:2778 PAD:13397 1.5
rPAD/9089 PAD:2778 PAD:13395 0.0375882
rPAD/9090 PAD:2778 PAD:13401 0.0751765
rPAD/9091 PAD:2754 PAD:13361 1.5
rPAD/9092 PAD:2754 PAD:13359 0.0375882
rPAD/9093 PAD:2754 PAD:13365 0.0751765
rPAD/9094 PAD:2750 PAD:13355 1.5
rPAD/9095 PAD:2750 PAD:13359 0.0751765
rPAD/9096 PAD:2748 PAD:13352 1.5
rPAD/9097 PAD:2748 PAD:2750 0.0375882
rPAD/9098 PAD:2746 PAD:13349 1.5
rPAD/9099 PAD:2746 PAD:13347 0.0375882
rPAD/9100 PAD:2746 PAD:2748 0.0751765
rPAD/9101 PAD:2742 PAD:13343 1.5
rPAD/9102 PAD:2742 PAD:13347 0.0751765
rPAD/9103 PAD:2740 PAD:13340 1.5
rPAD/9104 PAD:2740 PAD:13338 0.0751765
rPAD/9105 PAD:2740 PAD:2742 0.0375882
rPAD/9106 PAD:2726 PAD:13319 1.5
rPAD/9107 PAD:2726 PAD:13317 0.0375882
rPAD/9108 PAD:2726 PAD:13323 0.0751765
rPAD/9109 PAD:2718 PAD:13307 1.5
rPAD/9110 PAD:2718 PAD:13311 0.0751765
rPAD/9111 PAD:2716 PAD:13304 1.5
rPAD/9112 PAD:2716 PAD:2718 0.0375882
rPAD/9113 PAD:2714 PAD:13301 1.5
rPAD/9114 PAD:2714 PAD:2716 0.0751765
rPAD/9115 PAD:2712 PAD:13298 1.5
rPAD/9116 PAD:2712 PAD:2714 0.0375882
rPAD/9117 PAD:2710 PAD:13295 1.5
rPAD/9118 PAD:2710 PAD:13293 0.0375882
rPAD/9119 PAD:2710 PAD:2712 0.0751765
rPAD/9120 PAD:2704 PAD:13286 1.5
rPAD/9121 PAD:2704 PAD:13284 0.0751765
rPAD/9122 PAD:2704 PAD:13290 0.0375882
rPAD/9123 PAD:2690 PAD:13265 1.5
rPAD/9124 PAD:2690 PAD:13263 0.0375882
rPAD/9125 PAD:2690 PAD:13269 0.0751765
rPAD/9126 PAD:2673 PAD:2786 0.000694987
rPAD/9127 PAD:2673 PAD:13407 1.5
rPAD/9128 PAD:2673 PAD:13404 1.5
rPAD/9129 PAD:2673 PAD:13401 1.5
rPAD/9130 PAD:2673 PAD:2778 1.5
rPAD/9131 PAD:2673 PAD:13395 1.5
rPAD/9132 PAD:2673 PAD:13392 1.5
rPAD/9133 PAD:2673 PAD:13389 1.5
rPAD/9134 PAD:2673 PAD:13386 1.5
rPAD/9135 PAD:2673 PAD:13383 1.5
rPAD/9136 PAD:2673 PAD:13380 1.5
rPAD/9137 PAD:2673 PAD:13377 1.5
rPAD/9138 PAD:2673 PAD:13374 1.5
rPAD/9139 PAD:2673 PAD:13371 1.5
rPAD/9140 PAD:2673 PAD:13368 1.5
rPAD/9141 PAD:2673 PAD:13365 1.5
rPAD/9142 PAD:2673 PAD:2754 1.5
rPAD/9143 PAD:2673 PAD:13359 1.5
rPAD/9144 PAD:2673 PAD:2750 1.5
rPAD/9145 PAD:2673 PAD:2748 1.5
rPAD/9146 PAD:2673 PAD:2746 1.5
rPAD/9147 PAD:2673 PAD:13347 1.5
rPAD/9148 PAD:2673 PAD:2742 1.5
rPAD/9149 PAD:2673 PAD:2740 1.5
rPAD/9150 PAD:2673 PAD:13338 1.5
rPAD/9151 PAD:2673 PAD:13335 1.5
rPAD/9152 PAD:2673 PAD:13332 1.5
rPAD/9153 PAD:2673 PAD:13329 1.5
rPAD/9154 PAD:2673 PAD:13326 1.5
rPAD/9155 PAD:2673 PAD:13323 1.5
rPAD/9156 PAD:2673 PAD:2726 1.5
rPAD/9157 PAD:2673 PAD:13317 1.5
rPAD/9158 PAD:2673 PAD:13314 1.5
rPAD/9159 PAD:2673 PAD:13311 1.5
rPAD/9160 PAD:2673 PAD:2718 1.5
rPAD/9161 PAD:2673 PAD:2716 1.5
rPAD/9162 PAD:2673 PAD:2714 1.5
rPAD/9163 PAD:2673 PAD:2712 1.5
rPAD/9164 PAD:2673 PAD:2710 1.5
rPAD/9165 PAD:2673 PAD:13293 1.5
rPAD/9166 PAD:2673 PAD:13290 1.5
rPAD/9167 PAD:2673 PAD:2704 1.5
rPAD/9168 PAD:2673 PAD:13284 1.5
rPAD/9169 PAD:2673 PAD:13281 1.5
rPAD/9170 PAD:2673 PAD:13278 1.5
rPAD/9171 PAD:2673 PAD:13275 1.5
rPAD/9172 PAD:2673 PAD:13272 1.5
rPAD/9173 PAD:2673 PAD:13269 1.5
rPAD/9174 PAD:2673 PAD:2690 1.5
rPAD/9175 PAD:2673 PAD:13263 1.5
rPAD/9176 PAD:2673 PAD:13260 1.5
rPAD/9177 PAD:2673 PAD:13257 1.5
rPAD/9178 PAD:2673 PAD:13254 1.5
rPAD/9179 PAD:2673 PAD:13251 1.5
rPAD/9180 PAD:2673 PAD:13248 1.5
rPAD/9181 PAD:2673 PAD:13245 1.5
rPAD/9182 PAD:2673 PAD:13242 1.5
rPAD/9183 PAD:2670 PAD:2673 0.000174512
rPAD/9184 PAD:2670 PAD:14948 0.9
rPAD/9185 PAD:2668 PAD:16368 0.0285101
rPAD/9186 PAD:2668 PAD:15101 0.346154
rPAD/9187 PAD:2668 PAD:16426 0.0198121
rPAD/9188 PAD:2667 PAD:2670 9.49101e-05
rPAD/9189 PAD:2667 PAD:2668 0.346154
rPAD/9190 PAD:2659 PAD:13227 1.5
rPAD/9191 PAD:2659 PAD:13225 0.0375882
rPAD/9192 PAD:2659 PAD:13231 0.0751765
rPAD/9193 PAD:2635 PAD:13191 1.5
rPAD/9194 PAD:2635 PAD:13189 0.0375882
rPAD/9195 PAD:2635 PAD:13195 0.0751765
rPAD/9196 PAD:2631 PAD:13185 1.5
rPAD/9197 PAD:2631 PAD:13189 0.0751765
rPAD/9198 PAD:2629 PAD:13182 1.5
rPAD/9199 PAD:2629 PAD:2631 0.0375882
rPAD/9200 PAD:2627 PAD:13179 1.5
rPAD/9201 PAD:2627 PAD:13177 0.0375882
rPAD/9202 PAD:2627 PAD:2629 0.0751765
rPAD/9203 PAD:2623 PAD:13173 1.5
rPAD/9204 PAD:2623 PAD:13177 0.0751765
rPAD/9205 PAD:2621 PAD:13170 1.5
rPAD/9206 PAD:2621 PAD:13168 0.0751765
rPAD/9207 PAD:2621 PAD:2623 0.0375882
rPAD/9208 PAD:2607 PAD:13149 1.5
rPAD/9209 PAD:2607 PAD:13147 0.0375882
rPAD/9210 PAD:2607 PAD:13153 0.0751765
rPAD/9211 PAD:2599 PAD:13137 1.5
rPAD/9212 PAD:2599 PAD:13141 0.0751765
rPAD/9213 PAD:2597 PAD:13134 1.5
rPAD/9214 PAD:2597 PAD:2599 0.0375882
rPAD/9215 PAD:2595 PAD:13131 1.5
rPAD/9216 PAD:2595 PAD:2597 0.0751765
rPAD/9217 PAD:2593 PAD:13128 1.5
rPAD/9218 PAD:2593 PAD:2595 0.0375882
rPAD/9219 PAD:2591 PAD:13125 1.5
rPAD/9220 PAD:2591 PAD:13123 0.0375882
rPAD/9221 PAD:2591 PAD:2593 0.0751765
rPAD/9222 PAD:2585 PAD:13116 1.5
rPAD/9223 PAD:2585 PAD:13114 0.0751765
rPAD/9224 PAD:2585 PAD:13120 0.0375882
rPAD/9225 PAD:2571 PAD:13095 1.5
rPAD/9226 PAD:2571 PAD:13093 0.0375882
rPAD/9227 PAD:2571 PAD:13099 0.0751765
rPAD/9228 PAD:2554 PAD:2667 0.000946039
rPAD/9229 PAD:2554 PAD:13237 1.5
rPAD/9230 PAD:2554 PAD:13234 1.5
rPAD/9231 PAD:2554 PAD:13231 1.5
rPAD/9232 PAD:2554 PAD:2659 1.5
rPAD/9233 PAD:2554 PAD:13225 1.5
rPAD/9234 PAD:2554 PAD:13222 1.5
rPAD/9235 PAD:2554 PAD:13219 1.5
rPAD/9236 PAD:2554 PAD:13216 1.5
rPAD/9237 PAD:2554 PAD:13213 1.5
rPAD/9238 PAD:2554 PAD:13210 1.5
rPAD/9239 PAD:2554 PAD:13207 1.5
rPAD/9240 PAD:2554 PAD:13204 1.5
rPAD/9241 PAD:2554 PAD:13201 1.5
rPAD/9242 PAD:2554 PAD:13198 1.5
rPAD/9243 PAD:2554 PAD:13195 1.5
rPAD/9244 PAD:2554 PAD:2635 1.5
rPAD/9245 PAD:2554 PAD:13189 1.5
rPAD/9246 PAD:2554 PAD:2631 1.5
rPAD/9247 PAD:2554 PAD:2629 1.5
rPAD/9248 PAD:2554 PAD:2627 1.5
rPAD/9249 PAD:2554 PAD:13177 1.5
rPAD/9250 PAD:2554 PAD:2623 1.5
rPAD/9251 PAD:2554 PAD:2621 1.5
rPAD/9252 PAD:2554 PAD:13168 1.5
rPAD/9253 PAD:2554 PAD:13165 1.5
rPAD/9254 PAD:2554 PAD:13162 1.5
rPAD/9255 PAD:2554 PAD:13159 1.5
rPAD/9256 PAD:2554 PAD:13156 1.5
rPAD/9257 PAD:2554 PAD:13153 1.5
rPAD/9258 PAD:2554 PAD:2607 1.5
rPAD/9259 PAD:2554 PAD:13147 1.5
rPAD/9260 PAD:2554 PAD:13144 1.5
rPAD/9261 PAD:2554 PAD:13141 1.5
rPAD/9262 PAD:2554 PAD:2599 1.5
rPAD/9263 PAD:2554 PAD:2597 1.5
rPAD/9264 PAD:2554 PAD:2595 1.5
rPAD/9265 PAD:2554 PAD:2593 1.5
rPAD/9266 PAD:2554 PAD:2591 1.5
rPAD/9267 PAD:2554 PAD:13123 1.5
rPAD/9268 PAD:2554 PAD:13120 1.5
rPAD/9269 PAD:2554 PAD:2585 1.5
rPAD/9270 PAD:2554 PAD:13114 1.5
rPAD/9271 PAD:2554 PAD:13111 1.5
rPAD/9272 PAD:2554 PAD:13108 1.5
rPAD/9273 PAD:2554 PAD:13105 1.5
rPAD/9274 PAD:2554 PAD:13102 1.5
rPAD/9275 PAD:2554 PAD:13099 1.5
rPAD/9276 PAD:2554 PAD:2571 1.5
rPAD/9277 PAD:2554 PAD:13093 1.5
rPAD/9278 PAD:2554 PAD:13090 1.5
rPAD/9279 PAD:2554 PAD:13087 1.5
rPAD/9280 PAD:2554 PAD:13084 1.5
rPAD/9281 PAD:2554 PAD:13081 1.5
rPAD/9282 PAD:2554 PAD:13078 1.5
rPAD/9283 PAD:2554 PAD:13075 1.5
rPAD/9284 PAD:2554 PAD:13072 1.5
rPAD/9285 PAD:2552 PAD:16310 0.0318926
rPAD/9286 PAD:2552 PAD:15097 0.346154
rPAD/9287 PAD:2552 PAD:16368 0.0164295
rPAD/9288 PAD:2551 PAD:2554 0.000192882
rPAD/9289 PAD:2551 PAD:2552 0.346154
rPAD/9290 PAD:2548 PAD:2551 7.04171e-05
rPAD/9291 PAD:2548 PAD:14943 0.9
rPAD/9292 PAD:2545 PAD:2548 0.000869499
rPAD/9293 PAD:2545 PAD:14939 0.9
rPAD/9294 PAD:2537 PAD:13057 1.5
rPAD/9295 PAD:2537 PAD:13055 0.0375882
rPAD/9296 PAD:2537 PAD:13061 0.0751765
rPAD/9297 PAD:2513 PAD:13021 1.5
rPAD/9298 PAD:2513 PAD:13019 0.0375882
rPAD/9299 PAD:2513 PAD:13025 0.0751765
rPAD/9300 PAD:2509 PAD:13015 1.5
rPAD/9301 PAD:2509 PAD:13019 0.0751765
rPAD/9302 PAD:2507 PAD:13012 1.5
rPAD/9303 PAD:2507 PAD:2509 0.0375882
rPAD/9304 PAD:2505 PAD:13009 1.5
rPAD/9305 PAD:2505 PAD:13007 0.0375882
rPAD/9306 PAD:2505 PAD:2507 0.0751765
rPAD/9307 PAD:2501 PAD:13003 1.5
rPAD/9308 PAD:2501 PAD:13007 0.0751765
rPAD/9309 PAD:2499 PAD:13000 1.5
rPAD/9310 PAD:2499 PAD:12998 0.0751765
rPAD/9311 PAD:2499 PAD:2501 0.0375882
rPAD/9312 PAD:2485 PAD:12979 1.5
rPAD/9313 PAD:2485 PAD:12977 0.0375882
rPAD/9314 PAD:2485 PAD:12983 0.0751765
rPAD/9315 PAD:2477 PAD:12967 1.5
rPAD/9316 PAD:2477 PAD:12971 0.0751765
rPAD/9317 PAD:2475 PAD:12964 1.5
rPAD/9318 PAD:2475 PAD:2477 0.0375882
rPAD/9319 PAD:2473 PAD:12961 1.5
rPAD/9320 PAD:2473 PAD:2475 0.0751765
rPAD/9321 PAD:2471 PAD:12958 1.5
rPAD/9322 PAD:2471 PAD:2473 0.0375882
rPAD/9323 PAD:2469 PAD:12955 1.5
rPAD/9324 PAD:2469 PAD:12953 0.0375882
rPAD/9325 PAD:2469 PAD:2471 0.0751765
rPAD/9326 PAD:2463 PAD:12946 1.5
rPAD/9327 PAD:2463 PAD:12944 0.0751765
rPAD/9328 PAD:2463 PAD:12950 0.0375882
rPAD/9329 PAD:2449 PAD:12925 1.5
rPAD/9330 PAD:2449 PAD:12923 0.0375882
rPAD/9331 PAD:2449 PAD:12929 0.0751765
rPAD/9332 PAD:2432 PAD:2545 8.26636e-05
rPAD/9333 PAD:2432 PAD:13067 1.5
rPAD/9334 PAD:2432 PAD:13064 1.5
rPAD/9335 PAD:2432 PAD:13061 1.5
rPAD/9336 PAD:2432 PAD:2537 1.5
rPAD/9337 PAD:2432 PAD:13055 1.5
rPAD/9338 PAD:2432 PAD:13052 1.5
rPAD/9339 PAD:2432 PAD:13049 1.5
rPAD/9340 PAD:2432 PAD:13046 1.5
rPAD/9341 PAD:2432 PAD:13043 1.5
rPAD/9342 PAD:2432 PAD:13040 1.5
rPAD/9343 PAD:2432 PAD:13037 1.5
rPAD/9344 PAD:2432 PAD:13034 1.5
rPAD/9345 PAD:2432 PAD:13031 1.5
rPAD/9346 PAD:2432 PAD:13028 1.5
rPAD/9347 PAD:2432 PAD:13025 1.5
rPAD/9348 PAD:2432 PAD:2513 1.5
rPAD/9349 PAD:2432 PAD:13019 1.5
rPAD/9350 PAD:2432 PAD:2509 1.5
rPAD/9351 PAD:2432 PAD:2507 1.5
rPAD/9352 PAD:2432 PAD:2505 1.5
rPAD/9353 PAD:2432 PAD:13007 1.5
rPAD/9354 PAD:2432 PAD:2501 1.5
rPAD/9355 PAD:2432 PAD:2499 1.5
rPAD/9356 PAD:2432 PAD:12998 1.5
rPAD/9357 PAD:2432 PAD:12995 1.5
rPAD/9358 PAD:2432 PAD:12992 1.5
rPAD/9359 PAD:2432 PAD:12989 1.5
rPAD/9360 PAD:2432 PAD:12986 1.5
rPAD/9361 PAD:2432 PAD:12983 1.5
rPAD/9362 PAD:2432 PAD:2485 1.5
rPAD/9363 PAD:2432 PAD:12977 1.5
rPAD/9364 PAD:2432 PAD:12974 1.5
rPAD/9365 PAD:2432 PAD:12971 1.5
rPAD/9366 PAD:2432 PAD:2477 1.5
rPAD/9367 PAD:2432 PAD:2475 1.5
rPAD/9368 PAD:2432 PAD:2473 1.5
rPAD/9369 PAD:2432 PAD:2471 1.5
rPAD/9370 PAD:2432 PAD:2469 1.5
rPAD/9371 PAD:2432 PAD:12953 1.5
rPAD/9372 PAD:2432 PAD:12950 1.5
rPAD/9373 PAD:2432 PAD:2463 1.5
rPAD/9374 PAD:2432 PAD:12944 1.5
rPAD/9375 PAD:2432 PAD:12941 1.5
rPAD/9376 PAD:2432 PAD:12938 1.5
rPAD/9377 PAD:2432 PAD:12935 1.5
rPAD/9378 PAD:2432 PAD:12932 1.5
rPAD/9379 PAD:2432 PAD:12929 1.5
rPAD/9380 PAD:2432 PAD:2449 1.5
rPAD/9381 PAD:2432 PAD:12923 1.5
rPAD/9382 PAD:2432 PAD:12920 1.5
rPAD/9383 PAD:2432 PAD:12917 1.5
rPAD/9384 PAD:2432 PAD:12914 1.5
rPAD/9385 PAD:2432 PAD:12911 1.5
rPAD/9386 PAD:2432 PAD:12908 1.5
rPAD/9387 PAD:2432 PAD:12905 1.5
rPAD/9388 PAD:2432 PAD:12902 1.5
rPAD/9389 PAD:2430 PAD:16252 0.0352752
rPAD/9390 PAD:2430 PAD:9400 0.346154
rPAD/9391 PAD:2430 PAD:16310 0.013047
rPAD/9392 PAD:2429 PAD:2432 0.000116341
rPAD/9393 PAD:2429 PAD:2430 0.346154
rPAD/9394 PAD:2426 PAD:2429 0.00110524
rPAD/9395 PAD:2426 PAD:14934 0.9
rPAD/9396 PAD:2426 PAD:12897 1.5
rPAD/9397 PAD:2426 PAD:12894 1.5
rPAD/9398 PAD:2426 PAD:12891 1.5
rPAD/9399 PAD:2426 PAD:12885 1.5
rPAD/9400 PAD:2426 PAD:12882 1.5
rPAD/9401 PAD:2426 PAD:12879 1.5
rPAD/9402 PAD:2426 PAD:12876 1.5
rPAD/9403 PAD:2426 PAD:12873 1.5
rPAD/9404 PAD:2426 PAD:12870 1.5
rPAD/9405 PAD:2426 PAD:12867 1.5
rPAD/9406 PAD:2426 PAD:12864 1.5
rPAD/9407 PAD:2426 PAD:12861 1.5
rPAD/9408 PAD:2426 PAD:12858 1.5
rPAD/9409 PAD:2426 PAD:12855 1.5
rPAD/9410 PAD:2426 PAD:12849 1.5
rPAD/9411 PAD:2426 PAD:12837 1.5
rPAD/9412 PAD:2426 PAD:12828 1.5
rPAD/9413 PAD:2426 PAD:12825 1.5
rPAD/9414 PAD:2426 PAD:12822 1.5
rPAD/9415 PAD:2426 PAD:12819 1.5
rPAD/9416 PAD:2426 PAD:12816 1.5
rPAD/9417 PAD:2426 PAD:12813 1.5
rPAD/9418 PAD:2426 PAD:12807 1.5
rPAD/9419 PAD:2426 PAD:12804 1.5
rPAD/9420 PAD:2426 PAD:12801 1.5
rPAD/9421 PAD:2426 PAD:12783 1.5
rPAD/9422 PAD:2426 PAD:12780 1.5
rPAD/9423 PAD:2426 PAD:12774 1.5
rPAD/9424 PAD:2426 PAD:12771 1.5
rPAD/9425 PAD:2426 PAD:12768 1.5
rPAD/9426 PAD:2426 PAD:12765 1.5
rPAD/9427 PAD:2426 PAD:12762 1.5
rPAD/9428 PAD:2426 PAD:12759 1.5
rPAD/9429 PAD:2426 PAD:12753 1.5
rPAD/9430 PAD:2426 PAD:12750 1.5
rPAD/9431 PAD:2426 PAD:12747 1.5
rPAD/9432 PAD:2426 PAD:12744 1.5
rPAD/9433 PAD:2426 PAD:12741 1.5
rPAD/9434 PAD:2426 PAD:12738 1.5
rPAD/9435 PAD:2426 PAD:12735 1.5
rPAD/9436 PAD:2426 PAD:12732 1.5
rPAD/9437 PAD:2418 PAD:12887 1.5
rPAD/9438 PAD:2418 PAD:12885 0.0375882
rPAD/9439 PAD:2418 PAD:2426 1.5
rPAD/9440 PAD:2418 PAD:12891 0.0751765
rPAD/9441 PAD:2394 PAD:12851 1.5
rPAD/9442 PAD:2394 PAD:12849 0.0375882
rPAD/9443 PAD:2394 PAD:2426 1.5
rPAD/9444 PAD:2394 PAD:12855 0.0751765
rPAD/9445 PAD:2390 PAD:12845 1.5
rPAD/9446 PAD:2390 PAD:2426 1.5
rPAD/9447 PAD:2390 PAD:12849 0.0751765
rPAD/9448 PAD:2388 PAD:12842 1.5
rPAD/9449 PAD:2388 PAD:2426 1.5
rPAD/9450 PAD:2388 PAD:2390 0.0375882
rPAD/9451 PAD:2386 PAD:12839 1.5
rPAD/9452 PAD:2386 PAD:12837 0.0375882
rPAD/9453 PAD:2386 PAD:2426 1.5
rPAD/9454 PAD:2386 PAD:2388 0.0751765
rPAD/9455 PAD:2382 PAD:12833 1.5
rPAD/9456 PAD:2382 PAD:2426 1.5
rPAD/9457 PAD:2382 PAD:12837 0.0751765
rPAD/9458 PAD:2380 PAD:12830 1.5
rPAD/9459 PAD:2380 PAD:12828 0.0751765
rPAD/9460 PAD:2380 PAD:2426 1.5
rPAD/9461 PAD:2380 PAD:2382 0.0375882
rPAD/9462 PAD:2366 PAD:12809 1.5
rPAD/9463 PAD:2366 PAD:12807 0.0375882
rPAD/9464 PAD:2366 PAD:2426 1.5
rPAD/9465 PAD:2366 PAD:12813 0.0751765
rPAD/9466 PAD:2358 PAD:12797 1.5
rPAD/9467 PAD:2358 PAD:2426 1.5
rPAD/9468 PAD:2358 PAD:12801 0.0751765
rPAD/9469 PAD:2356 PAD:12794 1.5
rPAD/9470 PAD:2356 PAD:2426 1.5
rPAD/9471 PAD:2356 PAD:2358 0.0375882
rPAD/9472 PAD:2354 PAD:12791 1.5
rPAD/9473 PAD:2354 PAD:2426 1.5
rPAD/9474 PAD:2354 PAD:2356 0.0751765
rPAD/9475 PAD:2352 PAD:12788 1.5
rPAD/9476 PAD:2352 PAD:2426 1.5
rPAD/9477 PAD:2352 PAD:2354 0.0375882
rPAD/9478 PAD:2350 PAD:12785 1.5
rPAD/9479 PAD:2350 PAD:12783 0.0375882
rPAD/9480 PAD:2350 PAD:2426 1.5
rPAD/9481 PAD:2350 PAD:2352 0.0751765
rPAD/9482 PAD:2344 PAD:12776 1.5
rPAD/9483 PAD:2344 PAD:12774 0.0751765
rPAD/9484 PAD:2344 PAD:2426 1.5
rPAD/9485 PAD:2344 PAD:12780 0.0375882
rPAD/9486 PAD:2330 PAD:12755 1.5
rPAD/9487 PAD:2330 PAD:12753 0.0375882
rPAD/9488 PAD:2330 PAD:2426 1.5
rPAD/9489 PAD:2330 PAD:12759 0.0751765
rPAD/9490 PAD:2310 PAD:2426 3.06161e-05
rPAD/9491 PAD:2310 PAD:15090 0.346154
rPAD/9492 PAD:2307 PAD:2310 0.000835821
rPAD/9493 PAD:2307 PAD:14930 0.9
rPAD/9494 PAD:2299 PAD:12717 1.5
rPAD/9495 PAD:2299 PAD:12715 0.0375882
rPAD/9496 PAD:2299 PAD:12721 0.0751765
rPAD/9497 PAD:2275 PAD:12681 1.5
rPAD/9498 PAD:2275 PAD:12679 0.0375882
rPAD/9499 PAD:2275 PAD:12685 0.0751765
rPAD/9500 PAD:2271 PAD:12675 1.5
rPAD/9501 PAD:2271 PAD:12679 0.0751765
rPAD/9502 PAD:2269 PAD:12672 1.5
rPAD/9503 PAD:2269 PAD:2271 0.0375882
rPAD/9504 PAD:2267 PAD:12669 1.5
rPAD/9505 PAD:2267 PAD:12667 0.0375882
rPAD/9506 PAD:2267 PAD:2269 0.0751765
rPAD/9507 PAD:2263 PAD:12663 1.5
rPAD/9508 PAD:2263 PAD:12667 0.0751765
rPAD/9509 PAD:2261 PAD:12660 1.5
rPAD/9510 PAD:2261 PAD:12658 0.0751765
rPAD/9511 PAD:2261 PAD:2263 0.0375882
rPAD/9512 PAD:2247 PAD:12639 1.5
rPAD/9513 PAD:2247 PAD:12637 0.0375882
rPAD/9514 PAD:2247 PAD:12643 0.0751765
rPAD/9515 PAD:2239 PAD:12627 1.5
rPAD/9516 PAD:2239 PAD:12631 0.0751765
rPAD/9517 PAD:2237 PAD:12624 1.5
rPAD/9518 PAD:2237 PAD:2239 0.0375882
rPAD/9519 PAD:2235 PAD:12621 1.5
rPAD/9520 PAD:2235 PAD:2237 0.0751765
rPAD/9521 PAD:2233 PAD:12618 1.5
rPAD/9522 PAD:2233 PAD:2235 0.0375882
rPAD/9523 PAD:2231 PAD:12615 1.5
rPAD/9524 PAD:2231 PAD:12613 0.0375882
rPAD/9525 PAD:2231 PAD:2233 0.0751765
rPAD/9526 PAD:2225 PAD:12606 1.5
rPAD/9527 PAD:2225 PAD:12604 0.0751765
rPAD/9528 PAD:2225 PAD:12610 0.0375882
rPAD/9529 PAD:2211 PAD:12585 1.5
rPAD/9530 PAD:2211 PAD:12583 0.0375882
rPAD/9531 PAD:2211 PAD:12589 0.0751765
rPAD/9532 PAD:2194 PAD:2307 0.000361271
rPAD/9533 PAD:2194 PAD:12727 1.5
rPAD/9534 PAD:2194 PAD:12724 1.5
rPAD/9535 PAD:2194 PAD:12721 1.5
rPAD/9536 PAD:2194 PAD:2299 1.5
rPAD/9537 PAD:2194 PAD:12715 1.5
rPAD/9538 PAD:2194 PAD:12712 1.5
rPAD/9539 PAD:2194 PAD:12709 1.5
rPAD/9540 PAD:2194 PAD:12706 1.5
rPAD/9541 PAD:2194 PAD:12703 1.5
rPAD/9542 PAD:2194 PAD:12700 1.5
rPAD/9543 PAD:2194 PAD:12697 1.5
rPAD/9544 PAD:2194 PAD:12694 1.5
rPAD/9545 PAD:2194 PAD:12691 1.5
rPAD/9546 PAD:2194 PAD:12688 1.5
rPAD/9547 PAD:2194 PAD:12685 1.5
rPAD/9548 PAD:2194 PAD:2275 1.5
rPAD/9549 PAD:2194 PAD:12679 1.5
rPAD/9550 PAD:2194 PAD:2271 1.5
rPAD/9551 PAD:2194 PAD:2269 1.5
rPAD/9552 PAD:2194 PAD:2267 1.5
rPAD/9553 PAD:2194 PAD:12667 1.5
rPAD/9554 PAD:2194 PAD:2263 1.5
rPAD/9555 PAD:2194 PAD:2261 1.5
rPAD/9556 PAD:2194 PAD:12658 1.5
rPAD/9557 PAD:2194 PAD:12655 1.5
rPAD/9558 PAD:2194 PAD:12652 1.5
rPAD/9559 PAD:2194 PAD:12649 1.5
rPAD/9560 PAD:2194 PAD:12646 1.5
rPAD/9561 PAD:2194 PAD:12643 1.5
rPAD/9562 PAD:2194 PAD:2247 1.5
rPAD/9563 PAD:2194 PAD:12637 1.5
rPAD/9564 PAD:2194 PAD:12634 1.5
rPAD/9565 PAD:2194 PAD:12631 1.5
rPAD/9566 PAD:2194 PAD:2239 1.5
rPAD/9567 PAD:2194 PAD:2237 1.5
rPAD/9568 PAD:2194 PAD:2235 1.5
rPAD/9569 PAD:2194 PAD:2233 1.5
rPAD/9570 PAD:2194 PAD:2231 1.5
rPAD/9571 PAD:2194 PAD:12613 1.5
rPAD/9572 PAD:2194 PAD:12610 1.5
rPAD/9573 PAD:2194 PAD:2225 1.5
rPAD/9574 PAD:2194 PAD:12604 1.5
rPAD/9575 PAD:2194 PAD:12601 1.5
rPAD/9576 PAD:2194 PAD:12598 1.5
rPAD/9577 PAD:2194 PAD:12595 1.5
rPAD/9578 PAD:2194 PAD:12592 1.5
rPAD/9579 PAD:2194 PAD:12589 1.5
rPAD/9580 PAD:2194 PAD:2211 1.5
rPAD/9581 PAD:2194 PAD:12583 1.5
rPAD/9582 PAD:2194 PAD:12580 1.5
rPAD/9583 PAD:2194 PAD:12577 1.5
rPAD/9584 PAD:2194 PAD:12574 1.5
rPAD/9585 PAD:2194 PAD:12571 1.5
rPAD/9586 PAD:2194 PAD:12568 1.5
rPAD/9587 PAD:2194 PAD:12565 1.5
rPAD/9588 PAD:2194 PAD:12562 1.5
rPAD/9589 PAD:2191 PAD:2194 0.00032147
rPAD/9590 PAD:2191 PAD:15086 0.346154
rPAD/9591 PAD:2188 PAD:2191 0.000621508
rPAD/9592 PAD:2188 PAD:14924 0.9
rPAD/9593 PAD:2180 PAD:12547 1.5
rPAD/9594 PAD:2180 PAD:12545 0.0375882
rPAD/9595 PAD:2180 PAD:12551 0.0751765
rPAD/9596 PAD:2156 PAD:12511 1.5
rPAD/9597 PAD:2156 PAD:12509 0.0375882
rPAD/9598 PAD:2156 PAD:12515 0.0751765
rPAD/9599 PAD:2152 PAD:12505 1.5
rPAD/9600 PAD:2152 PAD:12509 0.0751765
rPAD/9601 PAD:2150 PAD:12502 1.5
rPAD/9602 PAD:2150 PAD:2152 0.0375882
rPAD/9603 PAD:2148 PAD:12499 1.5
rPAD/9604 PAD:2148 PAD:12497 0.0375882
rPAD/9605 PAD:2148 PAD:2150 0.0751765
rPAD/9606 PAD:2144 PAD:12493 1.5
rPAD/9607 PAD:2144 PAD:12497 0.0751765
rPAD/9608 PAD:2142 PAD:12490 1.5
rPAD/9609 PAD:2142 PAD:12488 0.0751765
rPAD/9610 PAD:2142 PAD:2144 0.0375882
rPAD/9611 PAD:2128 PAD:12469 1.5
rPAD/9612 PAD:2128 PAD:12467 0.0375882
rPAD/9613 PAD:2128 PAD:12473 0.0751765
rPAD/9614 PAD:2120 PAD:12457 1.5
rPAD/9615 PAD:2120 PAD:12461 0.0751765
rPAD/9616 PAD:2118 PAD:12454 1.5
rPAD/9617 PAD:2118 PAD:2120 0.0375882
rPAD/9618 PAD:2116 PAD:12451 1.5
rPAD/9619 PAD:2116 PAD:2118 0.0751765
rPAD/9620 PAD:2114 PAD:12448 1.5
rPAD/9621 PAD:2114 PAD:2116 0.0375882
rPAD/9622 PAD:2112 PAD:12445 1.5
rPAD/9623 PAD:2112 PAD:12443 0.0375882
rPAD/9624 PAD:2112 PAD:2114 0.0751765
rPAD/9625 PAD:2106 PAD:12436 1.5
rPAD/9626 PAD:2106 PAD:12434 0.0751765
rPAD/9627 PAD:2106 PAD:12440 0.0375882
rPAD/9628 PAD:2092 PAD:12415 1.5
rPAD/9629 PAD:2092 PAD:12413 0.0375882
rPAD/9630 PAD:2092 PAD:12419 0.0751765
rPAD/9631 PAD:2075 PAD:2188 0.000263299
rPAD/9632 PAD:2075 PAD:12557 1.5
rPAD/9633 PAD:2075 PAD:12554 1.5
rPAD/9634 PAD:2075 PAD:12551 1.5
rPAD/9635 PAD:2075 PAD:2180 1.5
rPAD/9636 PAD:2075 PAD:12545 1.5
rPAD/9637 PAD:2075 PAD:12542 1.5
rPAD/9638 PAD:2075 PAD:12539 1.5
rPAD/9639 PAD:2075 PAD:12536 1.5
rPAD/9640 PAD:2075 PAD:12533 1.5
rPAD/9641 PAD:2075 PAD:12530 1.5
rPAD/9642 PAD:2075 PAD:12527 1.5
rPAD/9643 PAD:2075 PAD:12524 1.5
rPAD/9644 PAD:2075 PAD:12521 1.5
rPAD/9645 PAD:2075 PAD:12518 1.5
rPAD/9646 PAD:2075 PAD:12515 1.5
rPAD/9647 PAD:2075 PAD:2156 1.5
rPAD/9648 PAD:2075 PAD:12509 1.5
rPAD/9649 PAD:2075 PAD:2152 1.5
rPAD/9650 PAD:2075 PAD:2150 1.5
rPAD/9651 PAD:2075 PAD:2148 1.5
rPAD/9652 PAD:2075 PAD:12497 1.5
rPAD/9653 PAD:2075 PAD:2144 1.5
rPAD/9654 PAD:2075 PAD:2142 1.5
rPAD/9655 PAD:2075 PAD:12488 1.5
rPAD/9656 PAD:2075 PAD:12485 1.5
rPAD/9657 PAD:2075 PAD:12482 1.5
rPAD/9658 PAD:2075 PAD:12479 1.5
rPAD/9659 PAD:2075 PAD:12476 1.5
rPAD/9660 PAD:2075 PAD:12473 1.5
rPAD/9661 PAD:2075 PAD:2128 1.5
rPAD/9662 PAD:2075 PAD:12467 1.5
rPAD/9663 PAD:2075 PAD:12464 1.5
rPAD/9664 PAD:2075 PAD:12461 1.5
rPAD/9665 PAD:2075 PAD:2120 1.5
rPAD/9666 PAD:2075 PAD:2118 1.5
rPAD/9667 PAD:2075 PAD:2116 1.5
rPAD/9668 PAD:2075 PAD:2114 1.5
rPAD/9669 PAD:2075 PAD:2112 1.5
rPAD/9670 PAD:2075 PAD:12443 1.5
rPAD/9671 PAD:2075 PAD:12440 1.5
rPAD/9672 PAD:2075 PAD:2106 1.5
rPAD/9673 PAD:2075 PAD:12434 1.5
rPAD/9674 PAD:2075 PAD:12431 1.5
rPAD/9675 PAD:2075 PAD:12428 1.5
rPAD/9676 PAD:2075 PAD:12425 1.5
rPAD/9677 PAD:2075 PAD:12422 1.5
rPAD/9678 PAD:2075 PAD:12419 1.5
rPAD/9679 PAD:2075 PAD:2092 1.5
rPAD/9680 PAD:2075 PAD:12413 1.5
rPAD/9681 PAD:2075 PAD:12410 1.5
rPAD/9682 PAD:2075 PAD:12407 1.5
rPAD/9683 PAD:2075 PAD:12404 1.5
rPAD/9684 PAD:2075 PAD:12401 1.5
rPAD/9685 PAD:2075 PAD:12398 1.5
rPAD/9686 PAD:2075 PAD:12395 1.5
rPAD/9687 PAD:2075 PAD:12392 1.5
rPAD/9688 PAD:2072 PAD:2075 0.000254114
rPAD/9689 PAD:2072 PAD:15082 0.346154
rPAD/9690 PAD:2070 PAD:16990 0.0269214
rPAD/9691 PAD:2070 PAD:9206 0.9
rPAD/9692 PAD:2070 PAD:16992 0.0516812
rPAD/9693 PAD:2069 PAD:2072 0.000352086
rPAD/9694 PAD:2069 PAD:2070 0.9
rPAD/9695 PAD:2061 PAD:12377 1.5
rPAD/9696 PAD:2061 PAD:12375 0.0375882
rPAD/9697 PAD:2061 PAD:12381 0.0751765
rPAD/9698 PAD:2037 PAD:12341 1.5
rPAD/9699 PAD:2037 PAD:12339 0.0375882
rPAD/9700 PAD:2037 PAD:12345 0.0751765
rPAD/9701 PAD:2033 PAD:12335 1.5
rPAD/9702 PAD:2033 PAD:12339 0.0751765
rPAD/9703 PAD:2031 PAD:12332 1.5
rPAD/9704 PAD:2031 PAD:2033 0.0375882
rPAD/9705 PAD:2029 PAD:12329 1.5
rPAD/9706 PAD:2029 PAD:12327 0.0375882
rPAD/9707 PAD:2029 PAD:2031 0.0751765
rPAD/9708 PAD:2025 PAD:12323 1.5
rPAD/9709 PAD:2025 PAD:12327 0.0751765
rPAD/9710 PAD:2023 PAD:12320 1.5
rPAD/9711 PAD:2023 PAD:12318 0.0751765
rPAD/9712 PAD:2023 PAD:2025 0.0375882
rPAD/9713 PAD:2009 PAD:12299 1.5
rPAD/9714 PAD:2009 PAD:12297 0.0375882
rPAD/9715 PAD:2009 PAD:12303 0.0751765
rPAD/9716 PAD:2001 PAD:12287 1.5
rPAD/9717 PAD:2001 PAD:12291 0.0751765
rPAD/9718 PAD:1999 PAD:12284 1.5
rPAD/9719 PAD:1999 PAD:2001 0.0375882
rPAD/9720 PAD:1997 PAD:12281 1.5
rPAD/9721 PAD:1997 PAD:1999 0.0751765
rPAD/9722 PAD:1995 PAD:12278 1.5
rPAD/9723 PAD:1995 PAD:1997 0.0375882
rPAD/9724 PAD:1993 PAD:12275 1.5
rPAD/9725 PAD:1993 PAD:12273 0.0375882
rPAD/9726 PAD:1993 PAD:1995 0.0751765
rPAD/9727 PAD:1987 PAD:12266 1.5
rPAD/9728 PAD:1987 PAD:12264 0.0751765
rPAD/9729 PAD:1987 PAD:12270 0.0375882
rPAD/9730 PAD:1973 PAD:12245 1.5
rPAD/9731 PAD:1973 PAD:12243 0.0375882
rPAD/9732 PAD:1973 PAD:12249 0.0751765
rPAD/9733 PAD:1956 PAD:2069 0.000627631
rPAD/9734 PAD:1956 PAD:12387 1.5
rPAD/9735 PAD:1956 PAD:12384 1.5
rPAD/9736 PAD:1956 PAD:12381 1.5
rPAD/9737 PAD:1956 PAD:2061 1.5
rPAD/9738 PAD:1956 PAD:12375 1.5
rPAD/9739 PAD:1956 PAD:12372 1.5
rPAD/9740 PAD:1956 PAD:12369 1.5
rPAD/9741 PAD:1956 PAD:12366 1.5
rPAD/9742 PAD:1956 PAD:12363 1.5
rPAD/9743 PAD:1956 PAD:12360 1.5
rPAD/9744 PAD:1956 PAD:12357 1.5
rPAD/9745 PAD:1956 PAD:12354 1.5
rPAD/9746 PAD:1956 PAD:12351 1.5
rPAD/9747 PAD:1956 PAD:12348 1.5
rPAD/9748 PAD:1956 PAD:12345 1.5
rPAD/9749 PAD:1956 PAD:2037 1.5
rPAD/9750 PAD:1956 PAD:12339 1.5
rPAD/9751 PAD:1956 PAD:2033 1.5
rPAD/9752 PAD:1956 PAD:2031 1.5
rPAD/9753 PAD:1956 PAD:2029 1.5
rPAD/9754 PAD:1956 PAD:12327 1.5
rPAD/9755 PAD:1956 PAD:2025 1.5
rPAD/9756 PAD:1956 PAD:2023 1.5
rPAD/9757 PAD:1956 PAD:12318 1.5
rPAD/9758 PAD:1956 PAD:12315 1.5
rPAD/9759 PAD:1956 PAD:12312 1.5
rPAD/9760 PAD:1956 PAD:12309 1.5
rPAD/9761 PAD:1956 PAD:12306 1.5
rPAD/9762 PAD:1956 PAD:12303 1.5
rPAD/9763 PAD:1956 PAD:2009 1.5
rPAD/9764 PAD:1956 PAD:12297 1.5
rPAD/9765 PAD:1956 PAD:12294 1.5
rPAD/9766 PAD:1956 PAD:12291 1.5
rPAD/9767 PAD:1956 PAD:2001 1.5
rPAD/9768 PAD:1956 PAD:1999 1.5
rPAD/9769 PAD:1956 PAD:1997 1.5
rPAD/9770 PAD:1956 PAD:1995 1.5
rPAD/9771 PAD:1956 PAD:1993 1.5
rPAD/9772 PAD:1956 PAD:12273 1.5
rPAD/9773 PAD:1956 PAD:12270 1.5
rPAD/9774 PAD:1956 PAD:1987 1.5
rPAD/9775 PAD:1956 PAD:12264 1.5
rPAD/9776 PAD:1956 PAD:12261 1.5
rPAD/9777 PAD:1956 PAD:12258 1.5
rPAD/9778 PAD:1956 PAD:12255 1.5
rPAD/9779 PAD:1956 PAD:12252 1.5
rPAD/9780 PAD:1956 PAD:12249 1.5
rPAD/9781 PAD:1956 PAD:1973 1.5
rPAD/9782 PAD:1956 PAD:12243 1.5
rPAD/9783 PAD:1956 PAD:12240 1.5
rPAD/9784 PAD:1956 PAD:12237 1.5
rPAD/9785 PAD:1956 PAD:12234 1.5
rPAD/9786 PAD:1956 PAD:12231 1.5
rPAD/9787 PAD:1956 PAD:12228 1.5
rPAD/9788 PAD:1956 PAD:12225 1.5
rPAD/9789 PAD:1956 PAD:12222 1.5
rPAD/9790 PAD:1954 PAD:16020 0.0338255
rPAD/9791 PAD:1954 PAD:9382 0.346154
rPAD/9792 PAD:1954 PAD:16078 0.0144966
rPAD/9793 PAD:1953 PAD:1956 0.000159204
rPAD/9794 PAD:1953 PAD:1954 0.346154
rPAD/9795 PAD:1951 PAD:16988 0.0218122
rPAD/9796 PAD:1951 PAD:14913 0.9
rPAD/9797 PAD:1951 PAD:16990 0.0567904
rPAD/9798 PAD:1950 PAD:1953 0.000517413
rPAD/9799 PAD:1950 PAD:1951 0.9
rPAD/9800 PAD PAD:1950 0.00039801
rPAD/9801 PAD:1940 PAD:12207 1.5
rPAD/9802 PAD:1940 PAD:12205 0.0375882
rPAD/9803 PAD:1940 PAD:12211 0.0751765
rPAD/9804 PAD:1916 PAD:12171 1.5
rPAD/9805 PAD:1916 PAD:12169 0.0375882
rPAD/9806 PAD:1916 PAD:12175 0.0751765
rPAD/9807 PAD:1912 PAD:12165 1.5
rPAD/9808 PAD:1912 PAD:12169 0.0751765
rPAD/9809 PAD:1910 PAD:12162 1.5
rPAD/9810 PAD:1910 PAD:1912 0.0375882
rPAD/9811 PAD:1908 PAD:12159 1.5
rPAD/9812 PAD:1908 PAD:12157 0.0375882
rPAD/9813 PAD:1908 PAD:1910 0.0751765
rPAD/9814 PAD:1904 PAD:12153 1.5
rPAD/9815 PAD:1904 PAD:12157 0.0751765
rPAD/9816 PAD:1902 PAD:12150 1.5
rPAD/9817 PAD:1902 PAD:12148 0.0751765
rPAD/9818 PAD:1902 PAD:1904 0.0375882
rPAD/9819 PAD:1888 PAD:12129 1.5
rPAD/9820 PAD:1888 PAD:12127 0.0375882
rPAD/9821 PAD:1888 PAD:12133 0.0751765
rPAD/9822 PAD:1880 PAD:12117 1.5
rPAD/9823 PAD:1880 PAD:12121 0.0751765
rPAD/9824 PAD:1878 PAD:12114 1.5
rPAD/9825 PAD:1878 PAD:1880 0.0375882
rPAD/9826 PAD:1876 PAD:12111 1.5
rPAD/9827 PAD:1876 PAD:1878 0.0751765
rPAD/9828 PAD:1874 PAD:12108 1.5
rPAD/9829 PAD:1874 PAD:1876 0.0375882
rPAD/9830 PAD:1872 PAD:12105 1.5
rPAD/9831 PAD:1872 PAD:12103 0.0375882
rPAD/9832 PAD:1872 PAD:1874 0.0751765
rPAD/9833 PAD:1866 PAD:12096 1.5
rPAD/9834 PAD:1866 PAD:12094 0.0751765
rPAD/9835 PAD:1866 PAD:12100 0.0375882
rPAD/9836 PAD:1852 PAD:12075 1.5
rPAD/9837 PAD:1852 PAD:12073 0.0375882
rPAD/9838 PAD:1852 PAD:12079 0.0751765
rPAD/9839 PAD:1835 PAD 0.000156142
rPAD/9840 PAD:1835 PAD:12217 1.5
rPAD/9841 PAD:1835 PAD:12214 1.5
rPAD/9842 PAD:1835 PAD:12211 1.5
rPAD/9843 PAD:1835 PAD:1940 1.5
rPAD/9844 PAD:1835 PAD:12205 1.5
rPAD/9845 PAD:1835 PAD:12202 1.5
rPAD/9846 PAD:1835 PAD:12199 1.5
rPAD/9847 PAD:1835 PAD:12196 1.5
rPAD/9848 PAD:1835 PAD:12193 1.5
rPAD/9849 PAD:1835 PAD:12190 1.5
rPAD/9850 PAD:1835 PAD:12187 1.5
rPAD/9851 PAD:1835 PAD:12184 1.5
rPAD/9852 PAD:1835 PAD:12181 1.5
rPAD/9853 PAD:1835 PAD:12178 1.5
rPAD/9854 PAD:1835 PAD:12175 1.5
rPAD/9855 PAD:1835 PAD:1916 1.5
rPAD/9856 PAD:1835 PAD:12169 1.5
rPAD/9857 PAD:1835 PAD:1912 1.5
rPAD/9858 PAD:1835 PAD:1910 1.5
rPAD/9859 PAD:1835 PAD:1908 1.5
rPAD/9860 PAD:1835 PAD:12157 1.5
rPAD/9861 PAD:1835 PAD:1904 1.5
rPAD/9862 PAD:1835 PAD:1902 1.5
rPAD/9863 PAD:1835 PAD:12148 1.5
rPAD/9864 PAD:1835 PAD:12145 1.5
rPAD/9865 PAD:1835 PAD:12142 1.5
rPAD/9866 PAD:1835 PAD:12139 1.5
rPAD/9867 PAD:1835 PAD:12136 1.5
rPAD/9868 PAD:1835 PAD:12133 1.5
rPAD/9869 PAD:1835 PAD:1888 1.5
rPAD/9870 PAD:1835 PAD:12127 1.5
rPAD/9871 PAD:1835 PAD:12124 1.5
rPAD/9872 PAD:1835 PAD:12121 1.5
rPAD/9873 PAD:1835 PAD:1880 1.5
rPAD/9874 PAD:1835 PAD:1878 1.5
rPAD/9875 PAD:1835 PAD:1876 1.5
rPAD/9876 PAD:1835 PAD:1874 1.5
rPAD/9877 PAD:1835 PAD:1872 1.5
rPAD/9878 PAD:1835 PAD:12103 1.5
rPAD/9879 PAD:1835 PAD:12100 1.5
rPAD/9880 PAD:1835 PAD:1866 1.5
rPAD/9881 PAD:1835 PAD:12094 1.5
rPAD/9882 PAD:1835 PAD:12091 1.5
rPAD/9883 PAD:1835 PAD:12088 1.5
rPAD/9884 PAD:1835 PAD:12085 1.5
rPAD/9885 PAD:1835 PAD:12082 1.5
rPAD/9886 PAD:1835 PAD:12079 1.5
rPAD/9887 PAD:1835 PAD:1852 1.5
rPAD/9888 PAD:1835 PAD:12073 1.5
rPAD/9889 PAD:1835 PAD:12070 1.5
rPAD/9890 PAD:1835 PAD:12067 1.5
rPAD/9891 PAD:1835 PAD:12064 1.5
rPAD/9892 PAD:1835 PAD:12061 1.5
rPAD/9893 PAD:1835 PAD:12058 1.5
rPAD/9894 PAD:1835 PAD:12055 1.5
rPAD/9895 PAD:1835 PAD:12052 1.5
rPAD/9896 PAD:1833 PAD:15962 0.0372081
rPAD/9897 PAD:1833 PAD:15073 0.346154
rPAD/9898 PAD:1833 PAD:16020 0.0111141
rPAD/9899 PAD:1832 PAD:1835 6.73555e-05
rPAD/9900 PAD:1832 PAD:1833 0.346154
rPAD/9901 PAD:1830 PAD:16986 0.044607
rPAD/9902 PAD:1830 PAD:14909 0.9
rPAD/9903 PAD:1830 PAD:16988 0.0339956
rPAD/9904 PAD:1829 PAD:1832 0.000247991
rPAD/9905 PAD:1829 PAD:1830 0.9
rPAD/9906 PAD:1821 PAD:12037 1.5
rPAD/9907 PAD:1821 PAD:12035 0.0375882
rPAD/9908 PAD:1821 PAD:12041 0.0751765
rPAD/9909 PAD:1797 PAD:12001 1.5
rPAD/9910 PAD:1797 PAD:11999 0.0375882
rPAD/9911 PAD:1797 PAD:12005 0.0751765
rPAD/9912 PAD:1793 PAD:11995 1.5
rPAD/9913 PAD:1793 PAD:11999 0.0751765
rPAD/9914 PAD:1791 PAD:11992 1.5
rPAD/9915 PAD:1791 PAD:1793 0.0375882
rPAD/9916 PAD:1789 PAD:11989 1.5
rPAD/9917 PAD:1789 PAD:11987 0.0375882
rPAD/9918 PAD:1789 PAD:1791 0.0751765
rPAD/9919 PAD:1785 PAD:11983 1.5
rPAD/9920 PAD:1785 PAD:11987 0.0751765
rPAD/9921 PAD:1783 PAD:11980 1.5
rPAD/9922 PAD:1783 PAD:11978 0.0751765
rPAD/9923 PAD:1783 PAD:1785 0.0375882
rPAD/9924 PAD:1769 PAD:11959 1.5
rPAD/9925 PAD:1769 PAD:11957 0.0375882
rPAD/9926 PAD:1769 PAD:11963 0.0751765
rPAD/9927 PAD:1761 PAD:11947 1.5
rPAD/9928 PAD:1761 PAD:11951 0.0751765
rPAD/9929 PAD:1759 PAD:11944 1.5
rPAD/9930 PAD:1759 PAD:1761 0.0375882
rPAD/9931 PAD:1757 PAD:11941 1.5
rPAD/9932 PAD:1757 PAD:1759 0.0751765
rPAD/9933 PAD:1755 PAD:11938 1.5
rPAD/9934 PAD:1755 PAD:1757 0.0375882
rPAD/9935 PAD:1753 PAD:11935 1.5
rPAD/9936 PAD:1753 PAD:11933 0.0375882
rPAD/9937 PAD:1753 PAD:1755 0.0751765
rPAD/9938 PAD:1747 PAD:11926 1.5
rPAD/9939 PAD:1747 PAD:11924 0.0751765
rPAD/9940 PAD:1747 PAD:11930 0.0375882
rPAD/9941 PAD:1733 PAD:11905 1.5
rPAD/9942 PAD:1733 PAD:11903 0.0375882
rPAD/9943 PAD:1733 PAD:11909 0.0751765
rPAD/9944 PAD:1716 PAD:1829 0.000918485
rPAD/9945 PAD:1716 PAD:12047 1.5
rPAD/9946 PAD:1716 PAD:12044 1.5
rPAD/9947 PAD:1716 PAD:12041 1.5
rPAD/9948 PAD:1716 PAD:1821 1.5
rPAD/9949 PAD:1716 PAD:12035 1.5
rPAD/9950 PAD:1716 PAD:12032 1.5
rPAD/9951 PAD:1716 PAD:12029 1.5
rPAD/9952 PAD:1716 PAD:12026 1.5
rPAD/9953 PAD:1716 PAD:12023 1.5
rPAD/9954 PAD:1716 PAD:12020 1.5
rPAD/9955 PAD:1716 PAD:12017 1.5
rPAD/9956 PAD:1716 PAD:12014 1.5
rPAD/9957 PAD:1716 PAD:12011 1.5
rPAD/9958 PAD:1716 PAD:12008 1.5
rPAD/9959 PAD:1716 PAD:12005 1.5
rPAD/9960 PAD:1716 PAD:1797 1.5
rPAD/9961 PAD:1716 PAD:11999 1.5
rPAD/9962 PAD:1716 PAD:1793 1.5
rPAD/9963 PAD:1716 PAD:1791 1.5
rPAD/9964 PAD:1716 PAD:1789 1.5
rPAD/9965 PAD:1716 PAD:11987 1.5
rPAD/9966 PAD:1716 PAD:1785 1.5
rPAD/9967 PAD:1716 PAD:1783 1.5
rPAD/9968 PAD:1716 PAD:11978 1.5
rPAD/9969 PAD:1716 PAD:11975 1.5
rPAD/9970 PAD:1716 PAD:11972 1.5
rPAD/9971 PAD:1716 PAD:11969 1.5
rPAD/9972 PAD:1716 PAD:11966 1.5
rPAD/9973 PAD:1716 PAD:11963 1.5
rPAD/9974 PAD:1716 PAD:1769 1.5
rPAD/9975 PAD:1716 PAD:11957 1.5
rPAD/9976 PAD:1716 PAD:11954 1.5
rPAD/9977 PAD:1716 PAD:11951 1.5
rPAD/9978 PAD:1716 PAD:1761 1.5
rPAD/9979 PAD:1716 PAD:1759 1.5
rPAD/9980 PAD:1716 PAD:1757 1.5
rPAD/9981 PAD:1716 PAD:1755 1.5
rPAD/9982 PAD:1716 PAD:1753 1.5
rPAD/9983 PAD:1716 PAD:11933 1.5
rPAD/9984 PAD:1716 PAD:11930 1.5
rPAD/9985 PAD:1716 PAD:1747 1.5
rPAD/9986 PAD:1716 PAD:11924 1.5
rPAD/9987 PAD:1716 PAD:11921 1.5
rPAD/9988 PAD:1716 PAD:11918 1.5
rPAD/9989 PAD:1716 PAD:11915 1.5
rPAD/9990 PAD:1716 PAD:11912 1.5
rPAD/9991 PAD:1716 PAD:11909 1.5
rPAD/9992 PAD:1716 PAD:1733 1.5
rPAD/9993 PAD:1716 PAD:11903 1.5
rPAD/9994 PAD:1716 PAD:11900 1.5
rPAD/9995 PAD:1716 PAD:11897 1.5
rPAD/9996 PAD:1716 PAD:11894 1.5
rPAD/9997 PAD:1716 PAD:11891 1.5
rPAD/9998 PAD:1716 PAD:11888 1.5
rPAD/9999 PAD:1716 PAD:11885 1.5
rPAD/10000 PAD:1716 PAD:11882 1.5
rPAD/10001 PAD:1714 PAD:15904 0.0256107
rPAD/10002 PAD:1714 PAD:15069 0.346154
rPAD/10003 PAD:1714 PAD:15962 0.0227114
rPAD/10004 PAD:1713 PAD:1716 0.000352086
rPAD/10005 PAD:1713 PAD:1714 0.346154
rPAD/10006 PAD:1711 PAD:16984 0.0394978
rPAD/10007 PAD:1711 PAD:14904 0.9
rPAD/10008 PAD:1711 PAD:16986 0.0391048
rPAD/10009 PAD:1710 PAD:1713 3.36778e-05
rPAD/10010 PAD:1710 PAD:1711 0.9
rPAD/10011 PAD:1702 PAD:11867 1.5
rPAD/10012 PAD:1702 PAD:11865 0.0375882
rPAD/10013 PAD:1702 PAD:11871 0.0751765
rPAD/10014 PAD:1678 PAD:11831 1.5
rPAD/10015 PAD:1678 PAD:11829 0.0375882
rPAD/10016 PAD:1678 PAD:11835 0.0751765
rPAD/10017 PAD:1674 PAD:11825 1.5
rPAD/10018 PAD:1674 PAD:11829 0.0751765
rPAD/10019 PAD:1672 PAD:11822 1.5
rPAD/10020 PAD:1672 PAD:1674 0.0375882
rPAD/10021 PAD:1670 PAD:11819 1.5
rPAD/10022 PAD:1670 PAD:11817 0.0375882
rPAD/10023 PAD:1670 PAD:1672 0.0751765
rPAD/10024 PAD:1666 PAD:11813 1.5
rPAD/10025 PAD:1666 PAD:11817 0.0751765
rPAD/10026 PAD:1664 PAD:11810 1.5
rPAD/10027 PAD:1664 PAD:11808 0.0751765
rPAD/10028 PAD:1664 PAD:1666 0.0375882
rPAD/10029 PAD:1650 PAD:11789 1.5
rPAD/10030 PAD:1650 PAD:11787 0.0375882
rPAD/10031 PAD:1650 PAD:11793 0.0751765
rPAD/10032 PAD:1642 PAD:11777 1.5
rPAD/10033 PAD:1642 PAD:11781 0.0751765
rPAD/10034 PAD:1640 PAD:11774 1.5
rPAD/10035 PAD:1640 PAD:1642 0.0375882
rPAD/10036 PAD:1638 PAD:11771 1.5
rPAD/10037 PAD:1638 PAD:1640 0.0751765
rPAD/10038 PAD:1636 PAD:11768 1.5
rPAD/10039 PAD:1636 PAD:1638 0.0375882
rPAD/10040 PAD:1634 PAD:11765 1.5
rPAD/10041 PAD:1634 PAD:11763 0.0375882
rPAD/10042 PAD:1634 PAD:1636 0.0751765
rPAD/10043 PAD:1628 PAD:11756 1.5
rPAD/10044 PAD:1628 PAD:11754 0.0751765
rPAD/10045 PAD:1628 PAD:11760 0.0375882
rPAD/10046 PAD:1614 PAD:11735 1.5
rPAD/10047 PAD:1614 PAD:11733 0.0375882
rPAD/10048 PAD:1614 PAD:11739 0.0751765
rPAD/10049 PAD:1597 PAD:1710 0.000829698
rPAD/10050 PAD:1597 PAD:11877 1.5
rPAD/10051 PAD:1597 PAD:11874 1.5
rPAD/10052 PAD:1597 PAD:11871 1.5
rPAD/10053 PAD:1597 PAD:1702 1.5
rPAD/10054 PAD:1597 PAD:11865 1.5
rPAD/10055 PAD:1597 PAD:11862 1.5
rPAD/10056 PAD:1597 PAD:11859 1.5
rPAD/10057 PAD:1597 PAD:11856 1.5
rPAD/10058 PAD:1597 PAD:11853 1.5
rPAD/10059 PAD:1597 PAD:11850 1.5
rPAD/10060 PAD:1597 PAD:11847 1.5
rPAD/10061 PAD:1597 PAD:11844 1.5
rPAD/10062 PAD:1597 PAD:11841 1.5
rPAD/10063 PAD:1597 PAD:11838 1.5
rPAD/10064 PAD:1597 PAD:11835 1.5
rPAD/10065 PAD:1597 PAD:1678 1.5
rPAD/10066 PAD:1597 PAD:11829 1.5
rPAD/10067 PAD:1597 PAD:1674 1.5
rPAD/10068 PAD:1597 PAD:1672 1.5
rPAD/10069 PAD:1597 PAD:1670 1.5
rPAD/10070 PAD:1597 PAD:11817 1.5
rPAD/10071 PAD:1597 PAD:1666 1.5
rPAD/10072 PAD:1597 PAD:1664 1.5
rPAD/10073 PAD:1597 PAD:11808 1.5
rPAD/10074 PAD:1597 PAD:11805 1.5
rPAD/10075 PAD:1597 PAD:11802 1.5
rPAD/10076 PAD:1597 PAD:11799 1.5
rPAD/10077 PAD:1597 PAD:11796 1.5
rPAD/10078 PAD:1597 PAD:11793 1.5
rPAD/10079 PAD:1597 PAD:1650 1.5
rPAD/10080 PAD:1597 PAD:11787 1.5
rPAD/10081 PAD:1597 PAD:11784 1.5
rPAD/10082 PAD:1597 PAD:11781 1.5
rPAD/10083 PAD:1597 PAD:1642 1.5
rPAD/10084 PAD:1597 PAD:1640 1.5
rPAD/10085 PAD:1597 PAD:1638 1.5
rPAD/10086 PAD:1597 PAD:1636 1.5
rPAD/10087 PAD:1597 PAD:1634 1.5
rPAD/10088 PAD:1597 PAD:11763 1.5
rPAD/10089 PAD:1597 PAD:11760 1.5
rPAD/10090 PAD:1597 PAD:1628 1.5
rPAD/10091 PAD:1597 PAD:11754 1.5
rPAD/10092 PAD:1597 PAD:11751 1.5
rPAD/10093 PAD:1597 PAD:11748 1.5
rPAD/10094 PAD:1597 PAD:11745 1.5
rPAD/10095 PAD:1597 PAD:11742 1.5
rPAD/10096 PAD:1597 PAD:11739 1.5
rPAD/10097 PAD:1597 PAD:1614 1.5
rPAD/10098 PAD:1597 PAD:11733 1.5
rPAD/10099 PAD:1597 PAD:11730 1.5
rPAD/10100 PAD:1597 PAD:11727 1.5
rPAD/10101 PAD:1597 PAD:11724 1.5
rPAD/10102 PAD:1597 PAD:11721 1.5
rPAD/10103 PAD:1597 PAD:11718 1.5
rPAD/10104 PAD:1597 PAD:11715 1.5
rPAD/10105 PAD:1597 PAD:11712 1.5
rPAD/10106 PAD:1595 PAD:16982 0.0622926
rPAD/10107 PAD:1595 PAD:14899 0.9
rPAD/10108 PAD:1595 PAD:16984 0.01631
rPAD/10109 PAD:1594 PAD:1597 3.9801e-05
rPAD/10110 PAD:1594 PAD:1595 0.9
rPAD/10111 PAD:1592 PAD:15846 0.0289933
rPAD/10112 PAD:1592 PAD:15065 0.346154
rPAD/10113 PAD:1592 PAD:15904 0.0193289
rPAD/10114 PAD:1591 PAD:1594 0.000235744
rPAD/10115 PAD:1591 PAD:1592 0.346154
rPAD/10116 PAD:1583 PAD:11697 1.5
rPAD/10117 PAD:1583 PAD:11695 0.0375882
rPAD/10118 PAD:1583 PAD:11701 0.0751765
rPAD/10119 PAD:1559 PAD:11661 1.5
rPAD/10120 PAD:1559 PAD:11659 0.0375882
rPAD/10121 PAD:1559 PAD:11665 0.0751765
rPAD/10122 PAD:1555 PAD:11655 1.5
rPAD/10123 PAD:1555 PAD:11659 0.0751765
rPAD/10124 PAD:1553 PAD:11652 1.5
rPAD/10125 PAD:1553 PAD:1555 0.0375882
rPAD/10126 PAD:1551 PAD:11649 1.5
rPAD/10127 PAD:1551 PAD:11647 0.0375882
rPAD/10128 PAD:1551 PAD:1553 0.0751765
rPAD/10129 PAD:1547 PAD:11643 1.5
rPAD/10130 PAD:1547 PAD:11647 0.0751765
rPAD/10131 PAD:1545 PAD:11640 1.5
rPAD/10132 PAD:1545 PAD:11638 0.0751765
rPAD/10133 PAD:1545 PAD:1547 0.0375882
rPAD/10134 PAD:1531 PAD:11619 1.5
rPAD/10135 PAD:1531 PAD:11617 0.0375882
rPAD/10136 PAD:1531 PAD:11623 0.0751765
rPAD/10137 PAD:1523 PAD:11607 1.5
rPAD/10138 PAD:1523 PAD:11611 0.0751765
rPAD/10139 PAD:1521 PAD:11604 1.5
rPAD/10140 PAD:1521 PAD:1523 0.0375882
rPAD/10141 PAD:1519 PAD:11601 1.5
rPAD/10142 PAD:1519 PAD:1521 0.0751765
rPAD/10143 PAD:1517 PAD:11598 1.5
rPAD/10144 PAD:1517 PAD:1519 0.0375882
rPAD/10145 PAD:1515 PAD:11595 1.5
rPAD/10146 PAD:1515 PAD:11593 0.0375882
rPAD/10147 PAD:1515 PAD:1517 0.0751765
rPAD/10148 PAD:1509 PAD:11586 1.5
rPAD/10149 PAD:1509 PAD:11584 0.0751765
rPAD/10150 PAD:1509 PAD:11590 0.0375882
rPAD/10151 PAD:1495 PAD:11565 1.5
rPAD/10152 PAD:1495 PAD:11563 0.0375882
rPAD/10153 PAD:1495 PAD:11569 0.0751765
rPAD/10154 PAD:1478 PAD:1591 0.000939916
rPAD/10155 PAD:1478 PAD:11707 1.5
rPAD/10156 PAD:1478 PAD:11704 1.5
rPAD/10157 PAD:1478 PAD:11701 1.5
rPAD/10158 PAD:1478 PAD:1583 1.5
rPAD/10159 PAD:1478 PAD:11695 1.5
rPAD/10160 PAD:1478 PAD:11692 1.5
rPAD/10161 PAD:1478 PAD:11689 1.5
rPAD/10162 PAD:1478 PAD:11686 1.5
rPAD/10163 PAD:1478 PAD:11683 1.5
rPAD/10164 PAD:1478 PAD:11680 1.5
rPAD/10165 PAD:1478 PAD:11677 1.5
rPAD/10166 PAD:1478 PAD:11674 1.5
rPAD/10167 PAD:1478 PAD:11671 1.5
rPAD/10168 PAD:1478 PAD:11668 1.5
rPAD/10169 PAD:1478 PAD:11665 1.5
rPAD/10170 PAD:1478 PAD:1559 1.5
rPAD/10171 PAD:1478 PAD:11659 1.5
rPAD/10172 PAD:1478 PAD:1555 1.5
rPAD/10173 PAD:1478 PAD:1553 1.5
rPAD/10174 PAD:1478 PAD:1551 1.5
rPAD/10175 PAD:1478 PAD:11647 1.5
rPAD/10176 PAD:1478 PAD:1547 1.5
rPAD/10177 PAD:1478 PAD:1545 1.5
rPAD/10178 PAD:1478 PAD:11638 1.5
rPAD/10179 PAD:1478 PAD:11635 1.5
rPAD/10180 PAD:1478 PAD:11632 1.5
rPAD/10181 PAD:1478 PAD:11629 1.5
rPAD/10182 PAD:1478 PAD:11626 1.5
rPAD/10183 PAD:1478 PAD:11623 1.5
rPAD/10184 PAD:1478 PAD:1531 1.5
rPAD/10185 PAD:1478 PAD:11617 1.5
rPAD/10186 PAD:1478 PAD:11614 1.5
rPAD/10187 PAD:1478 PAD:11611 1.5
rPAD/10188 PAD:1478 PAD:1523 1.5
rPAD/10189 PAD:1478 PAD:1521 1.5
rPAD/10190 PAD:1478 PAD:1519 1.5
rPAD/10191 PAD:1478 PAD:1517 1.5
rPAD/10192 PAD:1478 PAD:1515 1.5
rPAD/10193 PAD:1478 PAD:11593 1.5
rPAD/10194 PAD:1478 PAD:11590 1.5
rPAD/10195 PAD:1478 PAD:1509 1.5
rPAD/10196 PAD:1478 PAD:11584 1.5
rPAD/10197 PAD:1478 PAD:11581 1.5
rPAD/10198 PAD:1478 PAD:11578 1.5
rPAD/10199 PAD:1478 PAD:11575 1.5
rPAD/10200 PAD:1478 PAD:11572 1.5
rPAD/10201 PAD:1478 PAD:11569 1.5
rPAD/10202 PAD:1478 PAD:1495 1.5
rPAD/10203 PAD:1478 PAD:11563 1.5
rPAD/10204 PAD:1478 PAD:11560 1.5
rPAD/10205 PAD:1478 PAD:11557 1.5
rPAD/10206 PAD:1478 PAD:11554 1.5
rPAD/10207 PAD:1478 PAD:11551 1.5
rPAD/10208 PAD:1478 PAD:11548 1.5
rPAD/10209 PAD:1478 PAD:11545 1.5
rPAD/10210 PAD:1478 PAD:11542 1.5
rPAD/10211 PAD:1476 PAD:14893 0.9
rPAD/10212 PAD:1476 PAD:14890 0.0558079
rPAD/10213 PAD:1476 PAD:16982 0.0214192
rPAD/10214 PAD:1475 PAD:1478 0.000128588
rPAD/10215 PAD:1475 PAD:1476 0.9
rPAD/10216 PAD:1473 PAD:15788 0.0323758
rPAD/10217 PAD:1473 PAD:15061 0.346154
rPAD/10218 PAD:1473 PAD:15846 0.0159463
rPAD/10219 PAD:1472 PAD:1475 7.04171e-05
rPAD/10220 PAD:1472 PAD:1473 0.346154
rPAD/10221 PAD:1469 PAD:1472 0.000799082
rPAD/10222 PAD:1469 PAD:14890 0.9
rPAD/10223 PAD:1461 PAD:11527 1.5
rPAD/10224 PAD:1461 PAD:11525 0.0375882
rPAD/10225 PAD:1461 PAD:11531 0.0751765
rPAD/10226 PAD:1437 PAD:11491 1.5
rPAD/10227 PAD:1437 PAD:11489 0.0375882
rPAD/10228 PAD:1437 PAD:11495 0.0751765
rPAD/10229 PAD:1433 PAD:11485 1.5
rPAD/10230 PAD:1433 PAD:11489 0.0751765
rPAD/10231 PAD:1431 PAD:11482 1.5
rPAD/10232 PAD:1431 PAD:1433 0.0375882
rPAD/10233 PAD:1429 PAD:11479 1.5
rPAD/10234 PAD:1429 PAD:11477 0.0375882
rPAD/10235 PAD:1429 PAD:1431 0.0751765
rPAD/10236 PAD:1425 PAD:11473 1.5
rPAD/10237 PAD:1425 PAD:11477 0.0751765
rPAD/10238 PAD:1423 PAD:11470 1.5
rPAD/10239 PAD:1423 PAD:11468 0.0751765
rPAD/10240 PAD:1423 PAD:1425 0.0375882
rPAD/10241 PAD:1409 PAD:11449 1.5
rPAD/10242 PAD:1409 PAD:11447 0.0375882
rPAD/10243 PAD:1409 PAD:11453 0.0751765
rPAD/10244 PAD:1401 PAD:11437 1.5
rPAD/10245 PAD:1401 PAD:11441 0.0751765
rPAD/10246 PAD:1399 PAD:11434 1.5
rPAD/10247 PAD:1399 PAD:1401 0.0375882
rPAD/10248 PAD:1397 PAD:11431 1.5
rPAD/10249 PAD:1397 PAD:1399 0.0751765
rPAD/10250 PAD:1395 PAD:11428 1.5
rPAD/10251 PAD:1395 PAD:1397 0.0375882
rPAD/10252 PAD:1393 PAD:11425 1.5
rPAD/10253 PAD:1393 PAD:11423 0.0375882
rPAD/10254 PAD:1393 PAD:1395 0.0751765
rPAD/10255 PAD:1387 PAD:11416 1.5
rPAD/10256 PAD:1387 PAD:11414 0.0751765
rPAD/10257 PAD:1387 PAD:11420 0.0375882
rPAD/10258 PAD:1373 PAD:11395 1.5
rPAD/10259 PAD:1373 PAD:11393 0.0375882
rPAD/10260 PAD:1373 PAD:11399 0.0751765
rPAD/10261 PAD:1356 PAD:1469 0.000241868
rPAD/10262 PAD:1356 PAD:11537 1.5
rPAD/10263 PAD:1356 PAD:11534 1.5
rPAD/10264 PAD:1356 PAD:11531 1.5
rPAD/10265 PAD:1356 PAD:1461 1.5
rPAD/10266 PAD:1356 PAD:11525 1.5
rPAD/10267 PAD:1356 PAD:11522 1.5
rPAD/10268 PAD:1356 PAD:11519 1.5
rPAD/10269 PAD:1356 PAD:11516 1.5
rPAD/10270 PAD:1356 PAD:11513 1.5
rPAD/10271 PAD:1356 PAD:11510 1.5
rPAD/10272 PAD:1356 PAD:11507 1.5
rPAD/10273 PAD:1356 PAD:11504 1.5
rPAD/10274 PAD:1356 PAD:11501 1.5
rPAD/10275 PAD:1356 PAD:11498 1.5
rPAD/10276 PAD:1356 PAD:11495 1.5
rPAD/10277 PAD:1356 PAD:1437 1.5
rPAD/10278 PAD:1356 PAD:11489 1.5
rPAD/10279 PAD:1356 PAD:1433 1.5
rPAD/10280 PAD:1356 PAD:1431 1.5
rPAD/10281 PAD:1356 PAD:1429 1.5
rPAD/10282 PAD:1356 PAD:11477 1.5
rPAD/10283 PAD:1356 PAD:1425 1.5
rPAD/10284 PAD:1356 PAD:1423 1.5
rPAD/10285 PAD:1356 PAD:11468 1.5
rPAD/10286 PAD:1356 PAD:11465 1.5
rPAD/10287 PAD:1356 PAD:11462 1.5
rPAD/10288 PAD:1356 PAD:11459 1.5
rPAD/10289 PAD:1356 PAD:11456 1.5
rPAD/10290 PAD:1356 PAD:11453 1.5
rPAD/10291 PAD:1356 PAD:1409 1.5
rPAD/10292 PAD:1356 PAD:11447 1.5
rPAD/10293 PAD:1356 PAD:11444 1.5
rPAD/10294 PAD:1356 PAD:11441 1.5
rPAD/10295 PAD:1356 PAD:1401 1.5
rPAD/10296 PAD:1356 PAD:1399 1.5
rPAD/10297 PAD:1356 PAD:1397 1.5
rPAD/10298 PAD:1356 PAD:1395 1.5
rPAD/10299 PAD:1356 PAD:1393 1.5
rPAD/10300 PAD:1356 PAD:11423 1.5
rPAD/10301 PAD:1356 PAD:11420 1.5
rPAD/10302 PAD:1356 PAD:1387 1.5
rPAD/10303 PAD:1356 PAD:11414 1.5
rPAD/10304 PAD:1356 PAD:11411 1.5
rPAD/10305 PAD:1356 PAD:11408 1.5
rPAD/10306 PAD:1356 PAD:11405 1.5
rPAD/10307 PAD:1356 PAD:11402 1.5
rPAD/10308 PAD:1356 PAD:11399 1.5
rPAD/10309 PAD:1356 PAD:1373 1.5
rPAD/10310 PAD:1356 PAD:11393 1.5
rPAD/10311 PAD:1356 PAD:11390 1.5
rPAD/10312 PAD:1356 PAD:11387 1.5
rPAD/10313 PAD:1356 PAD:11384 1.5
rPAD/10314 PAD:1356 PAD:11381 1.5
rPAD/10315 PAD:1356 PAD:11378 1.5
rPAD/10316 PAD:1356 PAD:11375 1.5
rPAD/10317 PAD:1356 PAD:11372 1.5
rPAD/10318 PAD:1354 PAD:15730 0.0357584
rPAD/10319 PAD:1354 PAD:15057 0.346154
rPAD/10320 PAD:1354 PAD:15788 0.0125638
rPAD/10321 PAD:1353 PAD:1356 9.79717e-05
rPAD/10322 PAD:1353 PAD:1354 0.346154
rPAD/10323 PAD:1350 PAD:1353 0.000964409
rPAD/10324 PAD:1350 PAD:14884 0.9
rPAD/10325 PAD:1342 PAD:11357 1.5
rPAD/10326 PAD:1342 PAD:11355 0.0375882
rPAD/10327 PAD:1342 PAD:11361 0.0751765
rPAD/10328 PAD:1318 PAD:11321 1.5
rPAD/10329 PAD:1318 PAD:11319 0.0375882
rPAD/10330 PAD:1318 PAD:11325 0.0751765
rPAD/10331 PAD:1314 PAD:11315 1.5
rPAD/10332 PAD:1314 PAD:11319 0.0751765
rPAD/10333 PAD:1312 PAD:11312 1.5
rPAD/10334 PAD:1312 PAD:1314 0.0375882
rPAD/10335 PAD:1310 PAD:11309 1.5
rPAD/10336 PAD:1310 PAD:11307 0.0375882
rPAD/10337 PAD:1310 PAD:1312 0.0751765
rPAD/10338 PAD:1306 PAD:11303 1.5
rPAD/10339 PAD:1306 PAD:11307 0.0751765
rPAD/10340 PAD:1304 PAD:11300 1.5
rPAD/10341 PAD:1304 PAD:11298 0.0751765
rPAD/10342 PAD:1304 PAD:1306 0.0375882
rPAD/10343 PAD:1290 PAD:11279 1.5
rPAD/10344 PAD:1290 PAD:11277 0.0375882
rPAD/10345 PAD:1290 PAD:11283 0.0751765
rPAD/10346 PAD:1282 PAD:11267 1.5
rPAD/10347 PAD:1282 PAD:11271 0.0751765
rPAD/10348 PAD:1280 PAD:11264 1.5
rPAD/10349 PAD:1280 PAD:1282 0.0375882
rPAD/10350 PAD:1278 PAD:11261 1.5
rPAD/10351 PAD:1278 PAD:1280 0.0751765
rPAD/10352 PAD:1276 PAD:11258 1.5
rPAD/10353 PAD:1276 PAD:1278 0.0375882
rPAD/10354 PAD:1274 PAD:11255 1.5
rPAD/10355 PAD:1274 PAD:11253 0.0375882
rPAD/10356 PAD:1274 PAD:1276 0.0751765
rPAD/10357 PAD:1268 PAD:11246 1.5
rPAD/10358 PAD:1268 PAD:11244 0.0751765
rPAD/10359 PAD:1268 PAD:11250 0.0375882
rPAD/10360 PAD:1254 PAD:11225 1.5
rPAD/10361 PAD:1254 PAD:11223 0.0375882
rPAD/10362 PAD:1254 PAD:11229 0.0751765
rPAD/10363 PAD:1237 PAD:1350 0.000162266
rPAD/10364 PAD:1237 PAD:11367 1.5
rPAD/10365 PAD:1237 PAD:11364 1.5
rPAD/10366 PAD:1237 PAD:11361 1.5
rPAD/10367 PAD:1237 PAD:1342 1.5
rPAD/10368 PAD:1237 PAD:11355 1.5
rPAD/10369 PAD:1237 PAD:11352 1.5
rPAD/10370 PAD:1237 PAD:11349 1.5
rPAD/10371 PAD:1237 PAD:11346 1.5
rPAD/10372 PAD:1237 PAD:11343 1.5
rPAD/10373 PAD:1237 PAD:11340 1.5
rPAD/10374 PAD:1237 PAD:11337 1.5
rPAD/10375 PAD:1237 PAD:11334 1.5
rPAD/10376 PAD:1237 PAD:11331 1.5
rPAD/10377 PAD:1237 PAD:11328 1.5
rPAD/10378 PAD:1237 PAD:11325 1.5
rPAD/10379 PAD:1237 PAD:1318 1.5
rPAD/10380 PAD:1237 PAD:11319 1.5
rPAD/10381 PAD:1237 PAD:1314 1.5
rPAD/10382 PAD:1237 PAD:1312 1.5
rPAD/10383 PAD:1237 PAD:1310 1.5
rPAD/10384 PAD:1237 PAD:11307 1.5
rPAD/10385 PAD:1237 PAD:1306 1.5
rPAD/10386 PAD:1237 PAD:1304 1.5
rPAD/10387 PAD:1237 PAD:11298 1.5
rPAD/10388 PAD:1237 PAD:11295 1.5
rPAD/10389 PAD:1237 PAD:11292 1.5
rPAD/10390 PAD:1237 PAD:11289 1.5
rPAD/10391 PAD:1237 PAD:11286 1.5
rPAD/10392 PAD:1237 PAD:11283 1.5
rPAD/10393 PAD:1237 PAD:1290 1.5
rPAD/10394 PAD:1237 PAD:11277 1.5
rPAD/10395 PAD:1237 PAD:11274 1.5
rPAD/10396 PAD:1237 PAD:11271 1.5
rPAD/10397 PAD:1237 PAD:1282 1.5
rPAD/10398 PAD:1237 PAD:1280 1.5
rPAD/10399 PAD:1237 PAD:1278 1.5
rPAD/10400 PAD:1237 PAD:1276 1.5
rPAD/10401 PAD:1237 PAD:1274 1.5
rPAD/10402 PAD:1237 PAD:11253 1.5
rPAD/10403 PAD:1237 PAD:11250 1.5
rPAD/10404 PAD:1237 PAD:1268 1.5
rPAD/10405 PAD:1237 PAD:11244 1.5
rPAD/10406 PAD:1237 PAD:11241 1.5
rPAD/10407 PAD:1237 PAD:11238 1.5
rPAD/10408 PAD:1237 PAD:11235 1.5
rPAD/10409 PAD:1237 PAD:11232 1.5
rPAD/10410 PAD:1237 PAD:11229 1.5
rPAD/10411 PAD:1237 PAD:1254 1.5
rPAD/10412 PAD:1237 PAD:11223 1.5
rPAD/10413 PAD:1237 PAD:11220 1.5
rPAD/10414 PAD:1237 PAD:11217 1.5
rPAD/10415 PAD:1237 PAD:11214 1.5
rPAD/10416 PAD:1237 PAD:11211 1.5
rPAD/10417 PAD:1237 PAD:11208 1.5
rPAD/10418 PAD:1237 PAD:11205 1.5
rPAD/10419 PAD:1237 PAD:11202 1.5
rPAD/10420 PAD:1235 PAD:15672 0.0241611
rPAD/10421 PAD:1235 PAD:15053 0.346154
rPAD/10422 PAD:1235 PAD:15730 0.0241611
rPAD/10423 PAD:1234 PAD:1237 0.000391887
rPAD/10424 PAD:1234 PAD:1235 0.346154
rPAD/10425 PAD:1232 PAD:16975 0.0190611
rPAD/10426 PAD:1232 PAD:14880 0.9
rPAD/10427 PAD:1232 PAD:14884 0.0558079
rPAD/10428 PAD:1231 PAD:1234 0.000315346
rPAD/10429 PAD:1231 PAD:1232 0.9
rPAD/10430 PAD:1223 PAD:11187 1.5
rPAD/10431 PAD:1223 PAD:11185 0.0375882
rPAD/10432 PAD:1223 PAD:11191 0.0751765
rPAD/10433 PAD:1199 PAD:11151 1.5
rPAD/10434 PAD:1199 PAD:11149 0.0375882
rPAD/10435 PAD:1199 PAD:11155 0.0751765
rPAD/10436 PAD:1195 PAD:11145 1.5
rPAD/10437 PAD:1195 PAD:11149 0.0751765
rPAD/10438 PAD:1193 PAD:11142 1.5
rPAD/10439 PAD:1193 PAD:1195 0.0375882
rPAD/10440 PAD:1191 PAD:11139 1.5
rPAD/10441 PAD:1191 PAD:11137 0.0375882
rPAD/10442 PAD:1191 PAD:1193 0.0751765
rPAD/10443 PAD:1187 PAD:11133 1.5
rPAD/10444 PAD:1187 PAD:11137 0.0751765
rPAD/10445 PAD:1185 PAD:11130 1.5
rPAD/10446 PAD:1185 PAD:11128 0.0751765
rPAD/10447 PAD:1185 PAD:1187 0.0375882
rPAD/10448 PAD:1171 PAD:11109 1.5
rPAD/10449 PAD:1171 PAD:11107 0.0375882
rPAD/10450 PAD:1171 PAD:11113 0.0751765
rPAD/10451 PAD:1163 PAD:11097 1.5
rPAD/10452 PAD:1163 PAD:11101 0.0751765
rPAD/10453 PAD:1161 PAD:11094 1.5
rPAD/10454 PAD:1161 PAD:1163 0.0375882
rPAD/10455 PAD:1159 PAD:11091 1.5
rPAD/10456 PAD:1159 PAD:1161 0.0751765
rPAD/10457 PAD:1157 PAD:11088 1.5
rPAD/10458 PAD:1157 PAD:1159 0.0375882
rPAD/10459 PAD:1155 PAD:11085 1.5
rPAD/10460 PAD:1155 PAD:11083 0.0375882
rPAD/10461 PAD:1155 PAD:1157 0.0751765
rPAD/10462 PAD:1149 PAD:11076 1.5
rPAD/10463 PAD:1149 PAD:11074 0.0751765
rPAD/10464 PAD:1149 PAD:11080 0.0375882
rPAD/10465 PAD:1135 PAD:11055 1.5
rPAD/10466 PAD:1135 PAD:11053 0.0375882
rPAD/10467 PAD:1135 PAD:11059 0.0751765
rPAD/10468 PAD:1118 PAD:1231 0.000532721
rPAD/10469 PAD:1118 PAD:11197 1.5
rPAD/10470 PAD:1118 PAD:11194 1.5
rPAD/10471 PAD:1118 PAD:11191 1.5
rPAD/10472 PAD:1118 PAD:1223 1.5
rPAD/10473 PAD:1118 PAD:11185 1.5
rPAD/10474 PAD:1118 PAD:11182 1.5
rPAD/10475 PAD:1118 PAD:11179 1.5
rPAD/10476 PAD:1118 PAD:11176 1.5
rPAD/10477 PAD:1118 PAD:11173 1.5
rPAD/10478 PAD:1118 PAD:11170 1.5
rPAD/10479 PAD:1118 PAD:11167 1.5
rPAD/10480 PAD:1118 PAD:11164 1.5
rPAD/10481 PAD:1118 PAD:11161 1.5
rPAD/10482 PAD:1118 PAD:11158 1.5
rPAD/10483 PAD:1118 PAD:11155 1.5
rPAD/10484 PAD:1118 PAD:1199 1.5
rPAD/10485 PAD:1118 PAD:11149 1.5
rPAD/10486 PAD:1118 PAD:1195 1.5
rPAD/10487 PAD:1118 PAD:1193 1.5
rPAD/10488 PAD:1118 PAD:1191 1.5
rPAD/10489 PAD:1118 PAD:11137 1.5
rPAD/10490 PAD:1118 PAD:1187 1.5
rPAD/10491 PAD:1118 PAD:1185 1.5
rPAD/10492 PAD:1118 PAD:11128 1.5
rPAD/10493 PAD:1118 PAD:11125 1.5
rPAD/10494 PAD:1118 PAD:11122 1.5
rPAD/10495 PAD:1118 PAD:11119 1.5
rPAD/10496 PAD:1118 PAD:11116 1.5
rPAD/10497 PAD:1118 PAD:11113 1.5
rPAD/10498 PAD:1118 PAD:1171 1.5
rPAD/10499 PAD:1118 PAD:11107 1.5
rPAD/10500 PAD:1118 PAD:11104 1.5
rPAD/10501 PAD:1118 PAD:11101 1.5
rPAD/10502 PAD:1118 PAD:1163 1.5
rPAD/10503 PAD:1118 PAD:1161 1.5
rPAD/10504 PAD:1118 PAD:1159 1.5
rPAD/10505 PAD:1118 PAD:1157 1.5
rPAD/10506 PAD:1118 PAD:1155 1.5
rPAD/10507 PAD:1118 PAD:11083 1.5
rPAD/10508 PAD:1118 PAD:11080 1.5
rPAD/10509 PAD:1118 PAD:1149 1.5
rPAD/10510 PAD:1118 PAD:11074 1.5
rPAD/10511 PAD:1118 PAD:11071 1.5
rPAD/10512 PAD:1118 PAD:11068 1.5
rPAD/10513 PAD:1118 PAD:11065 1.5
rPAD/10514 PAD:1118 PAD:11062 1.5
rPAD/10515 PAD:1118 PAD:11059 1.5
rPAD/10516 PAD:1118 PAD:1135 1.5
rPAD/10517 PAD:1118 PAD:11053 1.5
rPAD/10518 PAD:1118 PAD:11050 1.5
rPAD/10519 PAD:1118 PAD:11047 1.5
rPAD/10520 PAD:1118 PAD:11044 1.5
rPAD/10521 PAD:1118 PAD:11041 1.5
rPAD/10522 PAD:1118 PAD:11038 1.5
rPAD/10523 PAD:1118 PAD:11035 1.5
rPAD/10524 PAD:1118 PAD:11032 1.5
rPAD/10525 PAD:1116 PAD:15614 0.0275436
rPAD/10526 PAD:1116 PAD:15049 0.346154
rPAD/10527 PAD:1116 PAD:15672 0.0207785
rPAD/10528 PAD:1115 PAD:1118 0.000290853
rPAD/10529 PAD:1115 PAD:1116 0.346154
rPAD/10530 PAD:1113 PAD:16973 0.013952
rPAD/10531 PAD:1113 PAD:14875 0.9
rPAD/10532 PAD:1113 PAD:16975 0.0646507
rPAD/10533 PAD:1112 PAD:1115 0.000480674
rPAD/10534 PAD:1112 PAD:1113 0.9
rPAD/10535 PAD:1104 PAD:11017 1.5
rPAD/10536 PAD:1104 PAD:11015 0.0375882
rPAD/10537 PAD:1104 PAD:11021 0.0751765
rPAD/10538 PAD:1080 PAD:10981 1.5
rPAD/10539 PAD:1080 PAD:10979 0.0375882
rPAD/10540 PAD:1080 PAD:10985 0.0751765
rPAD/10541 PAD:1076 PAD:10975 1.5
rPAD/10542 PAD:1076 PAD:10979 0.0751765
rPAD/10543 PAD:1074 PAD:10972 1.5
rPAD/10544 PAD:1074 PAD:1076 0.0375882
rPAD/10545 PAD:1072 PAD:10969 1.5
rPAD/10546 PAD:1072 PAD:10967 0.0375882
rPAD/10547 PAD:1072 PAD:1074 0.0751765
rPAD/10548 PAD:1068 PAD:10963 1.5
rPAD/10549 PAD:1068 PAD:10967 0.0751765
rPAD/10550 PAD:1066 PAD:10960 1.5
rPAD/10551 PAD:1066 PAD:10958 0.0751765
rPAD/10552 PAD:1066 PAD:1068 0.0375882
rPAD/10553 PAD:1052 PAD:10939 1.5
rPAD/10554 PAD:1052 PAD:10937 0.0375882
rPAD/10555 PAD:1052 PAD:10943 0.0751765
rPAD/10556 PAD:1044 PAD:10927 1.5
rPAD/10557 PAD:1044 PAD:10931 0.0751765
rPAD/10558 PAD:1042 PAD:10924 1.5
rPAD/10559 PAD:1042 PAD:1044 0.0375882
rPAD/10560 PAD:1040 PAD:10921 1.5
rPAD/10561 PAD:1040 PAD:1042 0.0751765
rPAD/10562 PAD:1038 PAD:10918 1.5
rPAD/10563 PAD:1038 PAD:1040 0.0375882
rPAD/10564 PAD:1036 PAD:10915 1.5
rPAD/10565 PAD:1036 PAD:10913 0.0375882
rPAD/10566 PAD:1036 PAD:1038 0.0751765
rPAD/10567 PAD:1030 PAD:10906 1.5
rPAD/10568 PAD:1030 PAD:10904 0.0751765
rPAD/10569 PAD:1030 PAD:10910 0.0375882
rPAD/10570 PAD:1016 PAD:10885 1.5
rPAD/10571 PAD:1016 PAD:10883 0.0375882
rPAD/10572 PAD:1016 PAD:10889 0.0751765
rPAD/10573 PAD:999 PAD:1112 0.000443934
rPAD/10574 PAD:999 PAD:11027 1.5
rPAD/10575 PAD:999 PAD:11024 1.5
rPAD/10576 PAD:999 PAD:11021 1.5
rPAD/10577 PAD:999 PAD:1104 1.5
rPAD/10578 PAD:999 PAD:11015 1.5
rPAD/10579 PAD:999 PAD:11012 1.5
rPAD/10580 PAD:999 PAD:11009 1.5
rPAD/10581 PAD:999 PAD:11006 1.5
rPAD/10582 PAD:999 PAD:11003 1.5
rPAD/10583 PAD:999 PAD:11000 1.5
rPAD/10584 PAD:999 PAD:10997 1.5
rPAD/10585 PAD:999 PAD:10994 1.5
rPAD/10586 PAD:999 PAD:10991 1.5
rPAD/10587 PAD:999 PAD:10988 1.5
rPAD/10588 PAD:999 PAD:10985 1.5
rPAD/10589 PAD:999 PAD:1080 1.5
rPAD/10590 PAD:999 PAD:10979 1.5
rPAD/10591 PAD:999 PAD:1076 1.5
rPAD/10592 PAD:999 PAD:1074 1.5
rPAD/10593 PAD:999 PAD:1072 1.5
rPAD/10594 PAD:999 PAD:10967 1.5
rPAD/10595 PAD:999 PAD:1068 1.5
rPAD/10596 PAD:999 PAD:1066 1.5
rPAD/10597 PAD:999 PAD:10958 1.5
rPAD/10598 PAD:999 PAD:10955 1.5
rPAD/10599 PAD:999 PAD:10952 1.5
rPAD/10600 PAD:999 PAD:10949 1.5
rPAD/10601 PAD:999 PAD:10946 1.5
rPAD/10602 PAD:999 PAD:10943 1.5
rPAD/10603 PAD:999 PAD:1052 1.5
rPAD/10604 PAD:999 PAD:10937 1.5
rPAD/10605 PAD:999 PAD:10934 1.5
rPAD/10606 PAD:999 PAD:10931 1.5
rPAD/10607 PAD:999 PAD:1044 1.5
rPAD/10608 PAD:999 PAD:1042 1.5
rPAD/10609 PAD:999 PAD:1040 1.5
rPAD/10610 PAD:999 PAD:1038 1.5
rPAD/10611 PAD:999 PAD:1036 1.5
rPAD/10612 PAD:999 PAD:10913 1.5
rPAD/10613 PAD:999 PAD:10910 1.5
rPAD/10614 PAD:999 PAD:1030 1.5
rPAD/10615 PAD:999 PAD:10904 1.5
rPAD/10616 PAD:999 PAD:10901 1.5
rPAD/10617 PAD:999 PAD:10898 1.5
rPAD/10618 PAD:999 PAD:10895 1.5
rPAD/10619 PAD:999 PAD:10892 1.5
rPAD/10620 PAD:999 PAD:10889 1.5
rPAD/10621 PAD:999 PAD:1016 1.5
rPAD/10622 PAD:999 PAD:10883 1.5
rPAD/10623 PAD:999 PAD:10880 1.5
rPAD/10624 PAD:999 PAD:10877 1.5
rPAD/10625 PAD:999 PAD:10874 1.5
rPAD/10626 PAD:999 PAD:10871 1.5
rPAD/10627 PAD:999 PAD:10868 1.5
rPAD/10628 PAD:999 PAD:10865 1.5
rPAD/10629 PAD:999 PAD:10862 1.5
rPAD/10630 PAD:997 PAD:15556 0.0309262
rPAD/10631 PAD:997 PAD:15045 0.346154
rPAD/10632 PAD:997 PAD:15614 0.017396
rPAD/10633 PAD:996 PAD:999 0.000214313
rPAD/10634 PAD:996 PAD:997 0.346154
rPAD/10635 PAD:994 PAD:16971 0.0367467
rPAD/10636 PAD:994 PAD:14870 0.9
rPAD/10637 PAD:994 PAD:16973 0.0418559
rPAD/10638 PAD:993 PAD:996 0.000211251
rPAD/10639 PAD:993 PAD:994 0.9
rPAD/10640 PAD:985 PAD:10847 1.5
rPAD/10641 PAD:985 PAD:10845 0.0375882
rPAD/10642 PAD:985 PAD:10851 0.0751765
rPAD/10643 PAD:961 PAD:10811 1.5
rPAD/10644 PAD:961 PAD:10809 0.0375882
rPAD/10645 PAD:961 PAD:10815 0.0751765
rPAD/10646 PAD:957 PAD:10805 1.5
rPAD/10647 PAD:957 PAD:10809 0.0751765
rPAD/10648 PAD:955 PAD:10802 1.5
rPAD/10649 PAD:955 PAD:957 0.0375882
rPAD/10650 PAD:953 PAD:10799 1.5
rPAD/10651 PAD:953 PAD:10797 0.0375882
rPAD/10652 PAD:953 PAD:955 0.0751765
rPAD/10653 PAD:949 PAD:10793 1.5
rPAD/10654 PAD:949 PAD:10797 0.0751765
rPAD/10655 PAD:947 PAD:10790 1.5
rPAD/10656 PAD:947 PAD:10788 0.0751765
rPAD/10657 PAD:947 PAD:949 0.0375882
rPAD/10658 PAD:933 PAD:10769 1.5
rPAD/10659 PAD:933 PAD:10767 0.0375882
rPAD/10660 PAD:933 PAD:10773 0.0751765
rPAD/10661 PAD:925 PAD:10757 1.5
rPAD/10662 PAD:925 PAD:10761 0.0751765
rPAD/10663 PAD:923 PAD:10754 1.5
rPAD/10664 PAD:923 PAD:925 0.0375882
rPAD/10665 PAD:921 PAD:10751 1.5
rPAD/10666 PAD:921 PAD:923 0.0751765
rPAD/10667 PAD:919 PAD:10748 1.5
rPAD/10668 PAD:919 PAD:921 0.0375882
rPAD/10669 PAD:917 PAD:10745 1.5
rPAD/10670 PAD:917 PAD:10743 0.0375882
rPAD/10671 PAD:917 PAD:919 0.0751765
rPAD/10672 PAD:911 PAD:10736 1.5
rPAD/10673 PAD:911 PAD:10734 0.0751765
rPAD/10674 PAD:911 PAD:10740 0.0375882
rPAD/10675 PAD:897 PAD:10715 1.5
rPAD/10676 PAD:897 PAD:10713 0.0375882
rPAD/10677 PAD:897 PAD:10719 0.0751765
rPAD/10678 PAD:880 PAD:993 0.000799082
rPAD/10679 PAD:880 PAD:10857 1.5
rPAD/10680 PAD:880 PAD:10854 1.5
rPAD/10681 PAD:880 PAD:10851 1.5
rPAD/10682 PAD:880 PAD:985 1.5
rPAD/10683 PAD:880 PAD:10845 1.5
rPAD/10684 PAD:880 PAD:10842 1.5
rPAD/10685 PAD:880 PAD:10839 1.5
rPAD/10686 PAD:880 PAD:10836 1.5
rPAD/10687 PAD:880 PAD:10833 1.5
rPAD/10688 PAD:880 PAD:10830 1.5
rPAD/10689 PAD:880 PAD:10827 1.5
rPAD/10690 PAD:880 PAD:10824 1.5
rPAD/10691 PAD:880 PAD:10821 1.5
rPAD/10692 PAD:880 PAD:10818 1.5
rPAD/10693 PAD:880 PAD:10815 1.5
rPAD/10694 PAD:880 PAD:961 1.5
rPAD/10695 PAD:880 PAD:10809 1.5
rPAD/10696 PAD:880 PAD:957 1.5
rPAD/10697 PAD:880 PAD:955 1.5
rPAD/10698 PAD:880 PAD:953 1.5
rPAD/10699 PAD:880 PAD:10797 1.5
rPAD/10700 PAD:880 PAD:949 1.5
rPAD/10701 PAD:880 PAD:947 1.5
rPAD/10702 PAD:880 PAD:10788 1.5
rPAD/10703 PAD:880 PAD:10785 1.5
rPAD/10704 PAD:880 PAD:10782 1.5
rPAD/10705 PAD:880 PAD:10779 1.5
rPAD/10706 PAD:880 PAD:10776 1.5
rPAD/10707 PAD:880 PAD:10773 1.5
rPAD/10708 PAD:880 PAD:933 1.5
rPAD/10709 PAD:880 PAD:10767 1.5
rPAD/10710 PAD:880 PAD:10764 1.5
rPAD/10711 PAD:880 PAD:10761 1.5
rPAD/10712 PAD:880 PAD:925 1.5
rPAD/10713 PAD:880 PAD:923 1.5
rPAD/10714 PAD:880 PAD:921 1.5
rPAD/10715 PAD:880 PAD:919 1.5
rPAD/10716 PAD:880 PAD:917 1.5
rPAD/10717 PAD:880 PAD:10743 1.5
rPAD/10718 PAD:880 PAD:10740 1.5
rPAD/10719 PAD:880 PAD:911 1.5
rPAD/10720 PAD:880 PAD:10734 1.5
rPAD/10721 PAD:880 PAD:10731 1.5
rPAD/10722 PAD:880 PAD:10728 1.5
rPAD/10723 PAD:880 PAD:10725 1.5
rPAD/10724 PAD:880 PAD:10722 1.5
rPAD/10725 PAD:880 PAD:10719 1.5
rPAD/10726 PAD:880 PAD:897 1.5
rPAD/10727 PAD:880 PAD:10713 1.5
rPAD/10728 PAD:880 PAD:10710 1.5
rPAD/10729 PAD:880 PAD:10707 1.5
rPAD/10730 PAD:880 PAD:10704 1.5
rPAD/10731 PAD:880 PAD:10701 1.5
rPAD/10732 PAD:880 PAD:10698 1.5
rPAD/10733 PAD:880 PAD:10695 1.5
rPAD/10734 PAD:880 PAD:10692 1.5
rPAD/10735 PAD:878 PAD:15498 0.0343087
rPAD/10736 PAD:878 PAD:9343 0.346154
rPAD/10737 PAD:878 PAD:15556 0.0140134
rPAD/10738 PAD:877 PAD:880 0.000128588
rPAD/10739 PAD:877 PAD:878 0.346154
rPAD/10740 PAD:874 PAD:877 0.000376579
rPAD/10741 PAD:874 PAD:14865 0.9
rPAD/10742 PAD:866 PAD:10677 1.5
rPAD/10743 PAD:866 PAD:10675 0.0375882
rPAD/10744 PAD:866 PAD:10681 0.0751765
rPAD/10745 PAD:842 PAD:10641 1.5
rPAD/10746 PAD:842 PAD:10639 0.0375882
rPAD/10747 PAD:842 PAD:10645 0.0751765
rPAD/10748 PAD:838 PAD:10635 1.5
rPAD/10749 PAD:838 PAD:10639 0.0751765
rPAD/10750 PAD:836 PAD:10632 1.5
rPAD/10751 PAD:836 PAD:838 0.0375882
rPAD/10752 PAD:834 PAD:10629 1.5
rPAD/10753 PAD:834 PAD:10627 0.0375882
rPAD/10754 PAD:834 PAD:836 0.0751765
rPAD/10755 PAD:830 PAD:10623 1.5
rPAD/10756 PAD:830 PAD:10627 0.0751765
rPAD/10757 PAD:828 PAD:10620 1.5
rPAD/10758 PAD:828 PAD:10618 0.0751765
rPAD/10759 PAD:828 PAD:830 0.0375882
rPAD/10760 PAD:814 PAD:10599 1.5
rPAD/10761 PAD:814 PAD:10597 0.0375882
rPAD/10762 PAD:814 PAD:10603 0.0751765
rPAD/10763 PAD:806 PAD:10587 1.5
rPAD/10764 PAD:806 PAD:10591 0.0751765
rPAD/10765 PAD:804 PAD:10584 1.5
rPAD/10766 PAD:804 PAD:806 0.0375882
rPAD/10767 PAD:802 PAD:10581 1.5
rPAD/10768 PAD:802 PAD:804 0.0751765
rPAD/10769 PAD:800 PAD:10578 1.5
rPAD/10770 PAD:800 PAD:802 0.0375882
rPAD/10771 PAD:798 PAD:10575 1.5
rPAD/10772 PAD:798 PAD:10573 0.0375882
rPAD/10773 PAD:798 PAD:800 0.0751765
rPAD/10774 PAD:792 PAD:10566 1.5
rPAD/10775 PAD:792 PAD:10564 0.0751765
rPAD/10776 PAD:792 PAD:10570 0.0375882
rPAD/10777 PAD:778 PAD:10545 1.5
rPAD/10778 PAD:778 PAD:10543 0.0375882
rPAD/10779 PAD:778 PAD:10549 0.0751765
rPAD/10780 PAD:761 PAD:874 0.000707233
rPAD/10781 PAD:761 PAD:10687 1.5
rPAD/10782 PAD:761 PAD:10684 1.5
rPAD/10783 PAD:761 PAD:10681 1.5
rPAD/10784 PAD:761 PAD:866 1.5
rPAD/10785 PAD:761 PAD:10675 1.5
rPAD/10786 PAD:761 PAD:10672 1.5
rPAD/10787 PAD:761 PAD:10669 1.5
rPAD/10788 PAD:761 PAD:10666 1.5
rPAD/10789 PAD:761 PAD:10663 1.5
rPAD/10790 PAD:761 PAD:10660 1.5
rPAD/10791 PAD:761 PAD:10657 1.5
rPAD/10792 PAD:761 PAD:10654 1.5
rPAD/10793 PAD:761 PAD:10651 1.5
rPAD/10794 PAD:761 PAD:10648 1.5
rPAD/10795 PAD:761 PAD:10645 1.5
rPAD/10796 PAD:761 PAD:842 1.5
rPAD/10797 PAD:761 PAD:10639 1.5
rPAD/10798 PAD:761 PAD:838 1.5
rPAD/10799 PAD:761 PAD:836 1.5
rPAD/10800 PAD:761 PAD:834 1.5
rPAD/10801 PAD:761 PAD:10627 1.5
rPAD/10802 PAD:761 PAD:830 1.5
rPAD/10803 PAD:761 PAD:828 1.5
rPAD/10804 PAD:761 PAD:10618 1.5
rPAD/10805 PAD:761 PAD:10615 1.5
rPAD/10806 PAD:761 PAD:10612 1.5
rPAD/10807 PAD:761 PAD:10609 1.5
rPAD/10808 PAD:761 PAD:10606 1.5
rPAD/10809 PAD:761 PAD:10603 1.5
rPAD/10810 PAD:761 PAD:814 1.5
rPAD/10811 PAD:761 PAD:10597 1.5
rPAD/10812 PAD:761 PAD:10594 1.5
rPAD/10813 PAD:761 PAD:10591 1.5
rPAD/10814 PAD:761 PAD:806 1.5
rPAD/10815 PAD:761 PAD:804 1.5
rPAD/10816 PAD:761 PAD:802 1.5
rPAD/10817 PAD:761 PAD:800 1.5
rPAD/10818 PAD:761 PAD:798 1.5
rPAD/10819 PAD:761 PAD:10573 1.5
rPAD/10820 PAD:761 PAD:10570 1.5
rPAD/10821 PAD:761 PAD:792 1.5
rPAD/10822 PAD:761 PAD:10564 1.5
rPAD/10823 PAD:761 PAD:10561 1.5
rPAD/10824 PAD:761 PAD:10558 1.5
rPAD/10825 PAD:761 PAD:10555 1.5
rPAD/10826 PAD:761 PAD:10552 1.5
rPAD/10827 PAD:761 PAD:10549 1.5
rPAD/10828 PAD:761 PAD:778 1.5
rPAD/10829 PAD:761 PAD:10543 1.5
rPAD/10830 PAD:761 PAD:10540 1.5
rPAD/10831 PAD:761 PAD:10537 1.5
rPAD/10832 PAD:761 PAD:10534 1.5
rPAD/10833 PAD:761 PAD:10531 1.5
rPAD/10834 PAD:761 PAD:10528 1.5
rPAD/10835 PAD:761 PAD:10525 1.5
rPAD/10836 PAD:761 PAD:10522 1.5
rPAD/10837 PAD:758 PAD:761 0.000162266
rPAD/10838 PAD:758 PAD:14860 0.9
rPAD/10839 PAD:755 PAD:758 0.000272484
rPAD/10840 PAD:755 PAD:15038 0.346154
rPAD/10841 PAD:747 PAD:10507 1.5
rPAD/10842 PAD:747 PAD:10505 0.0375882
rPAD/10843 PAD:747 PAD:10511 0.0751765
rPAD/10844 PAD:723 PAD:10471 1.5
rPAD/10845 PAD:723 PAD:10469 0.0375882
rPAD/10846 PAD:723 PAD:10475 0.0751765
rPAD/10847 PAD:719 PAD:10465 1.5
rPAD/10848 PAD:719 PAD:10469 0.0751765
rPAD/10849 PAD:717 PAD:10462 1.5
rPAD/10850 PAD:717 PAD:719 0.0375882
rPAD/10851 PAD:715 PAD:10459 1.5
rPAD/10852 PAD:715 PAD:10457 0.0375882
rPAD/10853 PAD:715 PAD:717 0.0751765
rPAD/10854 PAD:711 PAD:10453 1.5
rPAD/10855 PAD:711 PAD:10457 0.0751765
rPAD/10856 PAD:709 PAD:10450 1.5
rPAD/10857 PAD:709 PAD:10448 0.0751765
rPAD/10858 PAD:709 PAD:711 0.0375882
rPAD/10859 PAD:695 PAD:10429 1.5
rPAD/10860 PAD:695 PAD:10427 0.0375882
rPAD/10861 PAD:695 PAD:10433 0.0751765
rPAD/10862 PAD:687 PAD:10417 1.5
rPAD/10863 PAD:687 PAD:10421 0.0751765
rPAD/10864 PAD:685 PAD:10414 1.5
rPAD/10865 PAD:685 PAD:687 0.0375882
rPAD/10866 PAD:683 PAD:10411 1.5
rPAD/10867 PAD:683 PAD:685 0.0751765
rPAD/10868 PAD:681 PAD:10408 1.5
rPAD/10869 PAD:681 PAD:683 0.0375882
rPAD/10870 PAD:679 PAD:10405 1.5
rPAD/10871 PAD:679 PAD:10403 0.0375882
rPAD/10872 PAD:679 PAD:681 0.0751765
rPAD/10873 PAD:673 PAD:10396 1.5
rPAD/10874 PAD:673 PAD:10394 0.0751765
rPAD/10875 PAD:673 PAD:10400 0.0375882
rPAD/10876 PAD:659 PAD:10375 1.5
rPAD/10877 PAD:659 PAD:10373 0.0375882
rPAD/10878 PAD:659 PAD:10379 0.0751765
rPAD/10879 PAD:642 PAD:755 0.000802143
rPAD/10880 PAD:642 PAD:10517 1.5
rPAD/10881 PAD:642 PAD:10514 1.5
rPAD/10882 PAD:642 PAD:10511 1.5
rPAD/10883 PAD:642 PAD:747 1.5
rPAD/10884 PAD:642 PAD:10505 1.5
rPAD/10885 PAD:642 PAD:10502 1.5
rPAD/10886 PAD:642 PAD:10499 1.5
rPAD/10887 PAD:642 PAD:10496 1.5
rPAD/10888 PAD:642 PAD:10493 1.5
rPAD/10889 PAD:642 PAD:10490 1.5
rPAD/10890 PAD:642 PAD:10487 1.5
rPAD/10891 PAD:642 PAD:10484 1.5
rPAD/10892 PAD:642 PAD:10481 1.5
rPAD/10893 PAD:642 PAD:10478 1.5
rPAD/10894 PAD:642 PAD:10475 1.5
rPAD/10895 PAD:642 PAD:723 1.5
rPAD/10896 PAD:642 PAD:10469 1.5
rPAD/10897 PAD:642 PAD:719 1.5
rPAD/10898 PAD:642 PAD:717 1.5
rPAD/10899 PAD:642 PAD:715 1.5
rPAD/10900 PAD:642 PAD:10457 1.5
rPAD/10901 PAD:642 PAD:711 1.5
rPAD/10902 PAD:642 PAD:709 1.5
rPAD/10903 PAD:642 PAD:10448 1.5
rPAD/10904 PAD:642 PAD:10445 1.5
rPAD/10905 PAD:642 PAD:10442 1.5
rPAD/10906 PAD:642 PAD:10439 1.5
rPAD/10907 PAD:642 PAD:10436 1.5
rPAD/10908 PAD:642 PAD:10433 1.5
rPAD/10909 PAD:642 PAD:695 1.5
rPAD/10910 PAD:642 PAD:10427 1.5
rPAD/10911 PAD:642 PAD:10424 1.5
rPAD/10912 PAD:642 PAD:10421 1.5
rPAD/10913 PAD:642 PAD:687 1.5
rPAD/10914 PAD:642 PAD:685 1.5
rPAD/10915 PAD:642 PAD:683 1.5
rPAD/10916 PAD:642 PAD:681 1.5
rPAD/10917 PAD:642 PAD:679 1.5
rPAD/10918 PAD:642 PAD:10403 1.5
rPAD/10919 PAD:642 PAD:10400 1.5
rPAD/10920 PAD:642 PAD:673 1.5
rPAD/10921 PAD:642 PAD:10394 1.5
rPAD/10922 PAD:642 PAD:10391 1.5
rPAD/10923 PAD:642 PAD:10388 1.5
rPAD/10924 PAD:642 PAD:10385 1.5
rPAD/10925 PAD:642 PAD:10382 1.5
rPAD/10926 PAD:642 PAD:10379 1.5
rPAD/10927 PAD:642 PAD:659 1.5
rPAD/10928 PAD:642 PAD:10373 1.5
rPAD/10929 PAD:642 PAD:10370 1.5
rPAD/10930 PAD:642 PAD:10367 1.5
rPAD/10931 PAD:642 PAD:10364 1.5
rPAD/10932 PAD:642 PAD:10361 1.5
rPAD/10933 PAD:642 PAD:10358 1.5
rPAD/10934 PAD:642 PAD:10355 1.5
rPAD/10935 PAD:642 PAD:10352 1.5
rPAD/10936 PAD:639 PAD:642 0.000229621
rPAD/10937 PAD:639 PAD:14855 0.9
rPAD/10938 PAD:636 PAD:639 0.000107157
rPAD/10939 PAD:636 PAD:15034 0.346154
rPAD/10940 PAD:634 PAD:16963 0.0721179
rPAD/10941 PAD:634 PAD:14850 0.9
rPAD/10942 PAD:634 PAD:16965 0.00648472
rPAD/10943 PAD:633 PAD:636 0.000762342
rPAD/10944 PAD:633 PAD:634 0.9
rPAD/10945 PAD:625 PAD:10337 1.5
rPAD/10946 PAD:625 PAD:10335 0.0375882
rPAD/10947 PAD:625 PAD:10341 0.0751765
rPAD/10948 PAD:601 PAD:10301 1.5
rPAD/10949 PAD:601 PAD:10299 0.0375882
rPAD/10950 PAD:601 PAD:10305 0.0751765
rPAD/10951 PAD:597 PAD:10295 1.5
rPAD/10952 PAD:597 PAD:10299 0.0751765
rPAD/10953 PAD:595 PAD:10292 1.5
rPAD/10954 PAD:595 PAD:597 0.0375882
rPAD/10955 PAD:593 PAD:10289 1.5
rPAD/10956 PAD:593 PAD:10287 0.0375882
rPAD/10957 PAD:593 PAD:595 0.0751765
rPAD/10958 PAD:589 PAD:10283 1.5
rPAD/10959 PAD:589 PAD:10287 0.0751765
rPAD/10960 PAD:587 PAD:10280 1.5
rPAD/10961 PAD:587 PAD:10278 0.0751765
rPAD/10962 PAD:587 PAD:589 0.0375882
rPAD/10963 PAD:573 PAD:10259 1.5
rPAD/10964 PAD:573 PAD:10257 0.0375882
rPAD/10965 PAD:573 PAD:10263 0.0751765
rPAD/10966 PAD:565 PAD:10247 1.5
rPAD/10967 PAD:565 PAD:10251 0.0751765
rPAD/10968 PAD:563 PAD:10244 1.5
rPAD/10969 PAD:563 PAD:565 0.0375882
rPAD/10970 PAD:561 PAD:10241 1.5
rPAD/10971 PAD:561 PAD:563 0.0751765
rPAD/10972 PAD:559 PAD:10238 1.5
rPAD/10973 PAD:559 PAD:561 0.0375882
rPAD/10974 PAD:557 PAD:10235 1.5
rPAD/10975 PAD:557 PAD:10233 0.0375882
rPAD/10976 PAD:557 PAD:559 0.0751765
rPAD/10977 PAD:551 PAD:10226 1.5
rPAD/10978 PAD:551 PAD:10224 0.0751765
rPAD/10979 PAD:551 PAD:10230 0.0375882
rPAD/10980 PAD:537 PAD:10205 1.5
rPAD/10981 PAD:537 PAD:10203 0.0375882
rPAD/10982 PAD:537 PAD:10209 0.0751765
rPAD/10983 PAD:520 PAD:633 0.000116341
rPAD/10984 PAD:520 PAD:10347 1.5
rPAD/10985 PAD:520 PAD:10344 1.5
rPAD/10986 PAD:520 PAD:10341 1.5
rPAD/10987 PAD:520 PAD:625 1.5
rPAD/10988 PAD:520 PAD:10335 1.5
rPAD/10989 PAD:520 PAD:10332 1.5
rPAD/10990 PAD:520 PAD:10329 1.5
rPAD/10991 PAD:520 PAD:10326 1.5
rPAD/10992 PAD:520 PAD:10323 1.5
rPAD/10993 PAD:520 PAD:10320 1.5
rPAD/10994 PAD:520 PAD:10317 1.5
rPAD/10995 PAD:520 PAD:10314 1.5
rPAD/10996 PAD:520 PAD:10311 1.5
rPAD/10997 PAD:520 PAD:10308 1.5
rPAD/10998 PAD:520 PAD:10305 1.5
rPAD/10999 PAD:520 PAD:601 1.5
rPAD/11000 PAD:520 PAD:10299 1.5
rPAD/11001 PAD:520 PAD:597 1.5
rPAD/11002 PAD:520 PAD:595 1.5
rPAD/11003 PAD:520 PAD:593 1.5
rPAD/11004 PAD:520 PAD:10287 1.5
rPAD/11005 PAD:520 PAD:589 1.5
rPAD/11006 PAD:520 PAD:587 1.5
rPAD/11007 PAD:520 PAD:10278 1.5
rPAD/11008 PAD:520 PAD:10275 1.5
rPAD/11009 PAD:520 PAD:10272 1.5
rPAD/11010 PAD:520 PAD:10269 1.5
rPAD/11011 PAD:520 PAD:10266 1.5
rPAD/11012 PAD:520 PAD:10263 1.5
rPAD/11013 PAD:520 PAD:573 1.5
rPAD/11014 PAD:520 PAD:10257 1.5
rPAD/11015 PAD:520 PAD:10254 1.5
rPAD/11016 PAD:520 PAD:10251 1.5
rPAD/11017 PAD:520 PAD:565 1.5
rPAD/11018 PAD:520 PAD:563 1.5
rPAD/11019 PAD:520 PAD:561 1.5
rPAD/11020 PAD:520 PAD:559 1.5
rPAD/11021 PAD:520 PAD:557 1.5
rPAD/11022 PAD:520 PAD:10233 1.5
rPAD/11023 PAD:520 PAD:10230 1.5
rPAD/11024 PAD:520 PAD:551 1.5
rPAD/11025 PAD:520 PAD:10224 1.5
rPAD/11026 PAD:520 PAD:10221 1.5
rPAD/11027 PAD:520 PAD:10218 1.5
rPAD/11028 PAD:520 PAD:10215 1.5
rPAD/11029 PAD:520 PAD:10212 1.5
rPAD/11030 PAD:520 PAD:10209 1.5
rPAD/11031 PAD:520 PAD:537 1.5
rPAD/11032 PAD:520 PAD:10203 1.5
rPAD/11033 PAD:520 PAD:10200 1.5
rPAD/11034 PAD:520 PAD:10197 1.5
rPAD/11035 PAD:520 PAD:10194 1.5
rPAD/11036 PAD:520 PAD:10191 1.5
rPAD/11037 PAD:520 PAD:10188 1.5
rPAD/11038 PAD:520 PAD:10185 1.5
rPAD/11039 PAD:520 PAD:10182 1.5
rPAD/11040 PAD:517 PAD:520 0.000260237
rPAD/11041 PAD:517 PAD:15030 0.346154
rPAD/11042 PAD:514 PAD:517 0.000927669
rPAD/11043 PAD:514 PAD:14846 0.9
rPAD/11044 PAD:506 PAD:10167 1.5
rPAD/11045 PAD:506 PAD:10165 0.0375882
rPAD/11046 PAD:506 PAD:10171 0.0751765
rPAD/11047 PAD:482 PAD:10131 1.5
rPAD/11048 PAD:482 PAD:10129 0.0375882
rPAD/11049 PAD:482 PAD:10135 0.0751765
rPAD/11050 PAD:478 PAD:10125 1.5
rPAD/11051 PAD:478 PAD:10129 0.0751765
rPAD/11052 PAD:476 PAD:10122 1.5
rPAD/11053 PAD:476 PAD:478 0.0375882
rPAD/11054 PAD:474 PAD:10119 1.5
rPAD/11055 PAD:474 PAD:10117 0.0375882
rPAD/11056 PAD:474 PAD:476 0.0751765
rPAD/11057 PAD:470 PAD:10113 1.5
rPAD/11058 PAD:470 PAD:10117 0.0751765
rPAD/11059 PAD:468 PAD:10110 1.5
rPAD/11060 PAD:468 PAD:10108 0.0751765
rPAD/11061 PAD:468 PAD:470 0.0375882
rPAD/11062 PAD:454 PAD:10089 1.5
rPAD/11063 PAD:454 PAD:10087 0.0375882
rPAD/11064 PAD:454 PAD:10093 0.0751765
rPAD/11065 PAD:446 PAD:10077 1.5
rPAD/11066 PAD:446 PAD:10081 0.0751765
rPAD/11067 PAD:444 PAD:10074 1.5
rPAD/11068 PAD:444 PAD:446 0.0375882
rPAD/11069 PAD:442 PAD:10071 1.5
rPAD/11070 PAD:442 PAD:444 0.0751765
rPAD/11071 PAD:440 PAD:10068 1.5
rPAD/11072 PAD:440 PAD:442 0.0375882
rPAD/11073 PAD:438 PAD:10065 1.5
rPAD/11074 PAD:438 PAD:10063 0.0375882
rPAD/11075 PAD:438 PAD:440 0.0751765
rPAD/11076 PAD:432 PAD:10056 1.5
rPAD/11077 PAD:432 PAD:10054 0.0751765
rPAD/11078 PAD:432 PAD:10060 0.0375882
rPAD/11079 PAD:418 PAD:10035 1.5
rPAD/11080 PAD:418 PAD:10033 0.0375882
rPAD/11081 PAD:418 PAD:10039 0.0751765
rPAD/11082 PAD:401 PAD:514 2.75545e-05
rPAD/11083 PAD:401 PAD:10177 1.5
rPAD/11084 PAD:401 PAD:10174 1.5
rPAD/11085 PAD:401 PAD:10171 1.5
rPAD/11086 PAD:401 PAD:506 1.5
rPAD/11087 PAD:401 PAD:10165 1.5
rPAD/11088 PAD:401 PAD:10162 1.5
rPAD/11089 PAD:401 PAD:10159 1.5
rPAD/11090 PAD:401 PAD:10156 1.5
rPAD/11091 PAD:401 PAD:10153 1.5
rPAD/11092 PAD:401 PAD:10150 1.5
rPAD/11093 PAD:401 PAD:10147 1.5
rPAD/11094 PAD:401 PAD:10144 1.5
rPAD/11095 PAD:401 PAD:10141 1.5
rPAD/11096 PAD:401 PAD:10138 1.5
rPAD/11097 PAD:401 PAD:10135 1.5
rPAD/11098 PAD:401 PAD:482 1.5
rPAD/11099 PAD:401 PAD:10129 1.5
rPAD/11100 PAD:401 PAD:478 1.5
rPAD/11101 PAD:401 PAD:476 1.5
rPAD/11102 PAD:401 PAD:474 1.5
rPAD/11103 PAD:401 PAD:10117 1.5
rPAD/11104 PAD:401 PAD:470 1.5
rPAD/11105 PAD:401 PAD:468 1.5
rPAD/11106 PAD:401 PAD:10108 1.5
rPAD/11107 PAD:401 PAD:10105 1.5
rPAD/11108 PAD:401 PAD:10102 1.5
rPAD/11109 PAD:401 PAD:10099 1.5
rPAD/11110 PAD:401 PAD:10096 1.5
rPAD/11111 PAD:401 PAD:10093 1.5
rPAD/11112 PAD:401 PAD:454 1.5
rPAD/11113 PAD:401 PAD:10087 1.5
rPAD/11114 PAD:401 PAD:10084 1.5
rPAD/11115 PAD:401 PAD:10081 1.5
rPAD/11116 PAD:401 PAD:446 1.5
rPAD/11117 PAD:401 PAD:444 1.5
rPAD/11118 PAD:401 PAD:442 1.5
rPAD/11119 PAD:401 PAD:440 1.5
rPAD/11120 PAD:401 PAD:438 1.5
rPAD/11121 PAD:401 PAD:10063 1.5
rPAD/11122 PAD:401 PAD:10060 1.5
rPAD/11123 PAD:401 PAD:432 1.5
rPAD/11124 PAD:401 PAD:10054 1.5
rPAD/11125 PAD:401 PAD:10051 1.5
rPAD/11126 PAD:401 PAD:10048 1.5
rPAD/11127 PAD:401 PAD:10045 1.5
rPAD/11128 PAD:401 PAD:10042 1.5
rPAD/11129 PAD:401 PAD:10039 1.5
rPAD/11130 PAD:401 PAD:418 1.5
rPAD/11131 PAD:401 PAD:10033 1.5
rPAD/11132 PAD:401 PAD:10030 1.5
rPAD/11133 PAD:401 PAD:10027 1.5
rPAD/11134 PAD:401 PAD:10024 1.5
rPAD/11135 PAD:401 PAD:10021 1.5
rPAD/11136 PAD:401 PAD:10018 1.5
rPAD/11137 PAD:401 PAD:10015 1.5
rPAD/11138 PAD:401 PAD:10012 1.5
rPAD/11139 PAD:398 PAD:401 0.000183697
rPAD/11140 PAD:398 PAD:15026 0.346154
rPAD/11141 PAD:395 PAD:398 0.000658247
rPAD/11142 PAD:395 PAD:14842 0.9
rPAD/11143 PAD:387 PAD:9997 1.5
rPAD/11144 PAD:387 PAD:9995 0.0375882
rPAD/11145 PAD:387 PAD:10001 0.0751765
rPAD/11146 PAD:363 PAD:9961 1.5
rPAD/11147 PAD:363 PAD:9959 0.0375882
rPAD/11148 PAD:363 PAD:9965 0.0751765
rPAD/11149 PAD:359 PAD:9955 1.5
rPAD/11150 PAD:359 PAD:9959 0.0751765
rPAD/11151 PAD:357 PAD:9952 1.5
rPAD/11152 PAD:357 PAD:359 0.0375882
rPAD/11153 PAD:355 PAD:9949 1.5
rPAD/11154 PAD:355 PAD:9947 0.0375882
rPAD/11155 PAD:355 PAD:357 0.0751765
rPAD/11156 PAD:351 PAD:9943 1.5
rPAD/11157 PAD:351 PAD:9947 0.0751765
rPAD/11158 PAD:349 PAD:9940 1.5
rPAD/11159 PAD:349 PAD:9938 0.0751765
rPAD/11160 PAD:349 PAD:351 0.0375882
rPAD/11161 PAD:335 PAD:9919 1.5
rPAD/11162 PAD:335 PAD:9917 0.0375882
rPAD/11163 PAD:335 PAD:9923 0.0751765
rPAD/11164 PAD:327 PAD:9907 1.5
rPAD/11165 PAD:327 PAD:9911 0.0751765
rPAD/11166 PAD:325 PAD:9904 1.5
rPAD/11167 PAD:325 PAD:327 0.0375882
rPAD/11168 PAD:323 PAD:9901 1.5
rPAD/11169 PAD:323 PAD:325 0.0751765
rPAD/11170 PAD:321 PAD:9898 1.5
rPAD/11171 PAD:321 PAD:323 0.0375882
rPAD/11172 PAD:319 PAD:9895 1.5
rPAD/11173 PAD:319 PAD:9893 0.0375882
rPAD/11174 PAD:319 PAD:321 0.0751765
rPAD/11175 PAD:313 PAD:9886 1.5
rPAD/11176 PAD:313 PAD:9884 0.0751765
rPAD/11177 PAD:313 PAD:9890 0.0375882
rPAD/11178 PAD:299 PAD:9865 1.5
rPAD/11179 PAD:299 PAD:9863 0.0375882
rPAD/11180 PAD:299 PAD:9869 0.0751765
rPAD/11181 PAD:282 PAD:395 0.000382702
rPAD/11182 PAD:282 PAD:10007 1.5
rPAD/11183 PAD:282 PAD:10004 1.5
rPAD/11184 PAD:282 PAD:10001 1.5
rPAD/11185 PAD:282 PAD:387 1.5
rPAD/11186 PAD:282 PAD:9995 1.5
rPAD/11187 PAD:282 PAD:9992 1.5
rPAD/11188 PAD:282 PAD:9989 1.5
rPAD/11189 PAD:282 PAD:9986 1.5
rPAD/11190 PAD:282 PAD:9983 1.5
rPAD/11191 PAD:282 PAD:9980 1.5
rPAD/11192 PAD:282 PAD:9977 1.5
rPAD/11193 PAD:282 PAD:9974 1.5
rPAD/11194 PAD:282 PAD:9971 1.5
rPAD/11195 PAD:282 PAD:9968 1.5
rPAD/11196 PAD:282 PAD:9965 1.5
rPAD/11197 PAD:282 PAD:363 1.5
rPAD/11198 PAD:282 PAD:9959 1.5
rPAD/11199 PAD:282 PAD:359 1.5
rPAD/11200 PAD:282 PAD:357 1.5
rPAD/11201 PAD:282 PAD:355 1.5
rPAD/11202 PAD:282 PAD:9947 1.5
rPAD/11203 PAD:282 PAD:351 1.5
rPAD/11204 PAD:282 PAD:349 1.5
rPAD/11205 PAD:282 PAD:9938 1.5
rPAD/11206 PAD:282 PAD:9935 1.5
rPAD/11207 PAD:282 PAD:9932 1.5
rPAD/11208 PAD:282 PAD:9929 1.5
rPAD/11209 PAD:282 PAD:9926 1.5
rPAD/11210 PAD:282 PAD:9923 1.5
rPAD/11211 PAD:282 PAD:335 1.5
rPAD/11212 PAD:282 PAD:9917 1.5
rPAD/11213 PAD:282 PAD:9914 1.5
rPAD/11214 PAD:282 PAD:9911 1.5
rPAD/11215 PAD:282 PAD:327 1.5
rPAD/11216 PAD:282 PAD:325 1.5
rPAD/11217 PAD:282 PAD:323 1.5
rPAD/11218 PAD:282 PAD:321 1.5
rPAD/11219 PAD:282 PAD:319 1.5
rPAD/11220 PAD:282 PAD:9893 1.5
rPAD/11221 PAD:282 PAD:9890 1.5
rPAD/11222 PAD:282 PAD:313 1.5
rPAD/11223 PAD:282 PAD:9884 1.5
rPAD/11224 PAD:282 PAD:9881 1.5
rPAD/11225 PAD:282 PAD:9878 1.5
rPAD/11226 PAD:282 PAD:9875 1.5
rPAD/11227 PAD:282 PAD:9872 1.5
rPAD/11228 PAD:282 PAD:9869 1.5
rPAD/11229 PAD:282 PAD:299 1.5
rPAD/11230 PAD:282 PAD:9863 1.5
rPAD/11231 PAD:282 PAD:9860 1.5
rPAD/11232 PAD:282 PAD:9857 1.5
rPAD/11233 PAD:282 PAD:9854 1.5
rPAD/11234 PAD:282 PAD:9851 1.5
rPAD/11235 PAD:282 PAD:9848 1.5
rPAD/11236 PAD:282 PAD:9845 1.5
rPAD/11237 PAD:282 PAD:9842 1.5
rPAD/11238 PAD:280 PAD:15208 0.0212617
rPAD/11239 PAD:280 PAD:15021 0.346154
rPAD/11240 PAD:280 PAD:15266 0.0270604
rPAD/11241 PAD:279 PAD:282 0.000477612
rPAD/11242 PAD:279 PAD:280 0.346154
rPAD/11243 PAD:276 PAD:279 0.000443934
rPAD/11244 PAD:276 PAD:14836 0.9
rPAD/11245 PAD:268 PAD:9827 1.5
rPAD/11246 PAD:268 PAD:9825 0.0375882
rPAD/11247 PAD:268 PAD:9831 0.0751765
rPAD/11248 PAD:244 PAD:9791 1.5
rPAD/11249 PAD:244 PAD:9789 0.0375882
rPAD/11250 PAD:244 PAD:9795 0.0751765
rPAD/11251 PAD:240 PAD:9785 1.5
rPAD/11252 PAD:240 PAD:9789 0.0751765
rPAD/11253 PAD:238 PAD:9782 1.5
rPAD/11254 PAD:238 PAD:240 0.0375882
rPAD/11255 PAD:236 PAD:9779 1.5
rPAD/11256 PAD:236 PAD:9777 0.0375882
rPAD/11257 PAD:236 PAD:238 0.0751765
rPAD/11258 PAD:232 PAD:9773 1.5
rPAD/11259 PAD:232 PAD:9777 0.0751765
rPAD/11260 PAD:230 PAD:9770 1.5
rPAD/11261 PAD:230 PAD:9768 0.0751765
rPAD/11262 PAD:230 PAD:232 0.0375882
rPAD/11263 PAD:216 PAD:9749 1.5
rPAD/11264 PAD:216 PAD:9747 0.0375882
rPAD/11265 PAD:216 PAD:9753 0.0751765
rPAD/11266 PAD:208 PAD:9737 1.5
rPAD/11267 PAD:208 PAD:9741 0.0751765
rPAD/11268 PAD:206 PAD:9734 1.5
rPAD/11269 PAD:206 PAD:208 0.0375882
rPAD/11270 PAD:204 PAD:9731 1.5
rPAD/11271 PAD:204 PAD:206 0.0751765
rPAD/11272 PAD:202 PAD:9728 1.5
rPAD/11273 PAD:202 PAD:204 0.0375882
rPAD/11274 PAD:200 PAD:9725 1.5
rPAD/11275 PAD:200 PAD:9723 0.0375882
rPAD/11276 PAD:200 PAD:202 0.0751765
rPAD/11277 PAD:194 PAD:9716 1.5
rPAD/11278 PAD:194 PAD:9714 0.0751765
rPAD/11279 PAD:194 PAD:9720 0.0375882
rPAD/11280 PAD:180 PAD:9695 1.5
rPAD/11281 PAD:180 PAD:9693 0.0375882
rPAD/11282 PAD:180 PAD:9699 0.0751765
rPAD/11283 PAD:163 PAD:276 0.000306161
rPAD/11284 PAD:163 PAD:9837 1.5
rPAD/11285 PAD:163 PAD:9834 1.5
rPAD/11286 PAD:163 PAD:9831 1.5
rPAD/11287 PAD:163 PAD:268 1.5
rPAD/11288 PAD:163 PAD:9825 1.5
rPAD/11289 PAD:163 PAD:9822 1.5
rPAD/11290 PAD:163 PAD:9819 1.5
rPAD/11291 PAD:163 PAD:9816 1.5
rPAD/11292 PAD:163 PAD:9813 1.5
rPAD/11293 PAD:163 PAD:9810 1.5
rPAD/11294 PAD:163 PAD:9807 1.5
rPAD/11295 PAD:163 PAD:9804 1.5
rPAD/11296 PAD:163 PAD:9801 1.5
rPAD/11297 PAD:163 PAD:9798 1.5
rPAD/11298 PAD:163 PAD:9795 1.5
rPAD/11299 PAD:163 PAD:244 1.5
rPAD/11300 PAD:163 PAD:9789 1.5
rPAD/11301 PAD:163 PAD:240 1.5
rPAD/11302 PAD:163 PAD:238 1.5
rPAD/11303 PAD:163 PAD:236 1.5
rPAD/11304 PAD:163 PAD:9777 1.5
rPAD/11305 PAD:163 PAD:232 1.5
rPAD/11306 PAD:163 PAD:230 1.5
rPAD/11307 PAD:163 PAD:9768 1.5
rPAD/11308 PAD:163 PAD:9765 1.5
rPAD/11309 PAD:163 PAD:9762 1.5
rPAD/11310 PAD:163 PAD:9759 1.5
rPAD/11311 PAD:163 PAD:9756 1.5
rPAD/11312 PAD:163 PAD:9753 1.5
rPAD/11313 PAD:163 PAD:216 1.5
rPAD/11314 PAD:163 PAD:9747 1.5
rPAD/11315 PAD:163 PAD:9744 1.5
rPAD/11316 PAD:163 PAD:9741 1.5
rPAD/11317 PAD:163 PAD:208 1.5
rPAD/11318 PAD:163 PAD:206 1.5
rPAD/11319 PAD:163 PAD:204 1.5
rPAD/11320 PAD:163 PAD:202 1.5
rPAD/11321 PAD:163 PAD:200 1.5
rPAD/11322 PAD:163 PAD:9723 1.5
rPAD/11323 PAD:163 PAD:9720 1.5
rPAD/11324 PAD:163 PAD:194 1.5
rPAD/11325 PAD:163 PAD:9714 1.5
rPAD/11326 PAD:163 PAD:9711 1.5
rPAD/11327 PAD:163 PAD:9708 1.5
rPAD/11328 PAD:163 PAD:9705 1.5
rPAD/11329 PAD:163 PAD:9702 1.5
rPAD/11330 PAD:163 PAD:9699 1.5
rPAD/11331 PAD:163 PAD:180 1.5
rPAD/11332 PAD:163 PAD:9693 1.5
rPAD/11333 PAD:163 PAD:9690 1.5
rPAD/11334 PAD:163 PAD:9687 1.5
rPAD/11335 PAD:163 PAD:9684 1.5
rPAD/11336 PAD:163 PAD:9681 1.5
rPAD/11337 PAD:163 PAD:9678 1.5
rPAD/11338 PAD:163 PAD:9675 1.5
rPAD/11339 PAD:163 PAD:9672 1.5
rPAD/11340 PAD:161 PAD:15017 0.346154
rPAD/11341 PAD:161 PAD:15208 0.0236779
rPAD/11342 PAD:160 PAD:163 0.000388825
rPAD/11343 PAD:160 PAD:161 0.346154
rPAD/11344 PAD:157 PAD:160 0.000174512
rPAD/11345 PAD:157 PAD:14831 0.9
rPAD/11346 PAD:155 PAD:15145 0.0326174
rPAD/11347 PAD:155 PAD:15014 0.346154
rPAD/11348 PAD:155 PAD:161 0.0449396
rPAD/11349 PAD:154 PAD:157 0.000964409
rPAD/11350 PAD:154 PAD:155 0.346154
rPAD/11351 PAD:150 PAD:9651 0.586956
rPAD/11352 PAD:148 PAD:9640 0.586956
rPAD/11353 PAD:148 PAD:9638 0.01395
rPAD/11354 PAD:148 PAD:9645 0.0279
rPAD/11355 PAD:144 PAD:9619 0.586956
rPAD/11356 PAD:144 PAD:9617 0.01395
rPAD/11357 PAD:136 PAD:9577 0.586956
rPAD/11358 PAD:136 PAD:9574 0.0279
rPAD/11359 PAD:134 PAD:9566 0.586956
rPAD/11360 PAD:134 PAD:9564 0.01395
rPAD/11361 PAD:132 PAD:3860 0.586956
rPAD/11362 PAD:124 PAD:9513 0.586956
rPAD/11363 PAD:124 PAD:9511 0.01395
rPAD/11364 PAD:122 PAD:9500 0.0279
rPAD/11365 PAD:122 PAD:3815 0.586956
rPAD/11366 PAD:120 PAD:9492 0.586956
rPAD/11367 PAD:118 PAD:9481 0.586956
rPAD/11368 PAD:118 PAD:9486 0.0279
rPAD/11369 PAD:114 PAD:9460 0.586956
rPAD/11370 PAD:114 PAD:9458 0.01395
rPAD/11371 PAD:114 PAD:9465 0.0279
rPAD/11372 PAD:113 PAD:154 9.79717e-05
rPAD/11373 PAD:113 PAD:9663 0.586956
rPAD/11374 PAD:113 PAD:150 0.586956
rPAD/11375 PAD:113 PAD:148 0.586956
rPAD/11376 PAD:113 PAD:9631 0.586956
rPAD/11377 PAD:113 PAD:144 0.586956
rPAD/11378 PAD:113 PAD:9610 0.586956
rPAD/11379 PAD:113 PAD:9599 0.586956
rPAD/11380 PAD:113 PAD:9588 0.586956
rPAD/11381 PAD:113 PAD:136 0.586956
rPAD/11382 PAD:113 PAD:134 0.586956
rPAD/11383 PAD:113 PAD:132 0.586956
rPAD/11384 PAD:113 PAD:9546 0.586956
rPAD/11385 PAD:113 PAD:9535 0.586956
rPAD/11386 PAD:113 PAD:9525 0.586956
rPAD/11387 PAD:113 PAD:124 0.586956
rPAD/11388 PAD:113 PAD:122 0.586956
rPAD/11389 PAD:113 PAD:120 0.586956
rPAD/11390 PAD:113 PAD:118 0.586956
rPAD/11391 PAD:113 PAD:9472 0.586956
rPAD/11392 PAD:113 PAD:114 0.586956
rPAD/11393 PAD:110 PAD:113 0.00037964
rPAD/11394 PAD:110 PAD:14827 0.9
rPAD/11395 PAD:106 PAD:9658 0.586956
rPAD/11396 PAD:106 PAD:9663 0.0279
rPAD/11397 PAD:104 PAD:9647 0.586956
rPAD/11398 PAD:104 PAD:9645 0.01395
rPAD/11399 PAD:104 PAD:150 0.0279
rPAD/11400 PAD:100 PAD:9626 0.586956
rPAD/11401 PAD:100 PAD:9631 0.0279
rPAD/11402 PAD:94 PAD:9594 0.586956
rPAD/11403 PAD:94 PAD:9599 0.0279
rPAD/11404 PAD:92 PAD:9584 0.586956
rPAD/11405 PAD:92 PAD:9588 0.01395
rPAD/11406 PAD:86 PAD:9552 0.586956
rPAD/11407 PAD:86 PAD:132 0.0279
rPAD/11408 PAD:82 PAD:9531 0.586956
rPAD/11409 PAD:82 PAD:9535 0.01395
rPAD/11410 PAD:80 PAD:9520 0.586956
rPAD/11411 PAD:80 PAD:9525 0.0279
rPAD/11412 PAD:74 PAD:9488 0.586956
rPAD/11413 PAD:74 PAD:9486 0.01395
rPAD/11414 PAD:74 PAD:120 0.0279
rPAD/11415 PAD:72 PAD:9478 0.586956
rPAD/11416 PAD:72 PAD:9476 0.01395
rPAD/11417 PAD:72 PAD:118 0.01395
rPAD/11418 PAD:70 PAD:9467 0.586956
rPAD/11419 PAD:70 PAD:9465 0.01395
rPAD/11420 PAD:70 PAD:9472 0.0279
rPAD/11421 PAD:65 PAD:110 0.00037964
rPAD/11422 PAD:65 PAD:9666 0.225
rPAD/11423 PAD:65 PAD:106 0.586956
rPAD/11424 PAD:65 PAD:104 0.586956
rPAD/11425 PAD:65 PAD:9638 0.586956
rPAD/11426 PAD:65 PAD:100 0.586956
rPAD/11427 PAD:65 PAD:9617 0.586956
rPAD/11428 PAD:65 PAD:9606 0.586956
rPAD/11429 PAD:65 PAD:94 0.586956
rPAD/11430 PAD:65 PAD:92 0.586956
rPAD/11431 PAD:65 PAD:9574 0.586956
rPAD/11432 PAD:65 PAD:9564 0.586956
rPAD/11433 PAD:65 PAD:86 0.586956
rPAD/11434 PAD:65 PAD:9542 0.586956
rPAD/11435 PAD:65 PAD:82 0.586956
rPAD/11436 PAD:65 PAD:80 0.586956
rPAD/11437 PAD:65 PAD:9511 0.586956
rPAD/11438 PAD:65 PAD:9500 0.586956
rPAD/11439 PAD:65 PAD:74 0.586956
rPAD/11440 PAD:65 PAD:72 0.586956
rPAD/11441 PAD:65 PAD:70 0.586956
rPAD/11442 PAD:65 PAD:9458 0.586956
rPAD/11443 PAD:65 PAD:14823 0.9
rPAD/11444 PAD:63 PAD:15008 0.346154
rPAD/11445 PAD:63 PAD:15145 0.0123221
rPAD/11446 PAD:62 PAD:65 0.000281669
rPAD/11447 PAD:62 PAD:63 0.346154
rPAD/11448 PAD:60 PAD:9655 0.586956
rPAD/11449 PAD:60 PAD:150 0.0279
rPAD/11450 PAD:60 PAD:106 0.01395
rPAD/11451 PAD:56 PAD:9634 0.586956
rPAD/11452 PAD:56 PAD:9631 0.0279
rPAD/11453 PAD:56 PAD:9638 0.01395
rPAD/11454 PAD:54 PAD:9623 0.586956
rPAD/11455 PAD:54 PAD:144 0.0279
rPAD/11456 PAD:54 PAD:100 0.01395
rPAD/11457 PAD:48 PAD:9591 0.586956
rPAD/11458 PAD:48 PAD:9588 0.0279
rPAD/11459 PAD:48 PAD:94 0.01395
rPAD/11460 PAD:46 PAD:9581 0.586956
rPAD/11461 PAD:46 PAD:136 0.0279
rPAD/11462 PAD:46 PAD:92 0.01395
rPAD/11463 PAD:44 PAD:9570 0.586956
rPAD/11464 PAD:44 PAD:134 0.0279
rPAD/11465 PAD:44 PAD:9574 0.01395
rPAD/11466 PAD:42 PAD:9559 0.586956
rPAD/11467 PAD:42 PAD:132 0.01395
rPAD/11468 PAD:42 PAD:9564 0.0279
rPAD/11469 PAD:40 PAD:9549 0.586956
rPAD/11470 PAD:40 PAD:9546 0.0279
rPAD/11471 PAD:40 PAD:86 0.01395
rPAD/11472 PAD:38 PAD:9538 0.586956
rPAD/11473 PAD:38 PAD:9535 0.0279
rPAD/11474 PAD:38 PAD:9542 0.01395
rPAD/11475 PAD:36 PAD:9528 0.586956
rPAD/11476 PAD:36 PAD:9525 0.0279
rPAD/11477 PAD:36 PAD:82 0.01395
rPAD/11478 PAD:34 PAD:9517 0.586956
rPAD/11479 PAD:34 PAD:124 0.0279
rPAD/11480 PAD:34 PAD:80 0.01395
rPAD/11481 PAD:32 PAD:9506 0.586956
rPAD/11482 PAD:32 PAD:122 0.01395
rPAD/11483 PAD:32 PAD:9511 0.0279
rPAD/11484 PAD:30 PAD:9496 0.586956
rPAD/11485 PAD:30 PAD:120 0.0279
rPAD/11486 PAD:30 PAD:9500 0.01395
rPAD/11487 PAD:19 PAD:9086 0.9
rPAD/11488 PAD:19 PAD:14823 0.0487336
rPAD/11489 PAD:18 PAD:62 0.000477612
rPAD/11490 PAD:18 PAD:60 0.586956
rPAD/11491 PAD:18 PAD:9645 0.586956
rPAD/11492 PAD:18 PAD:56 0.586956
rPAD/11493 PAD:18 PAD:54 0.586956
rPAD/11494 PAD:18 PAD:9613 0.586956
rPAD/11495 PAD:18 PAD:9603 0.586956
rPAD/11496 PAD:18 PAD:48 0.586956
rPAD/11497 PAD:18 PAD:46 0.586956
rPAD/11498 PAD:18 PAD:44 0.586956
rPAD/11499 PAD:18 PAD:42 0.586956
rPAD/11500 PAD:18 PAD:40 0.586956
rPAD/11501 PAD:18 PAD:38 0.586956
rPAD/11502 PAD:18 PAD:36 0.586956
rPAD/11503 PAD:18 PAD:34 0.586956
rPAD/11504 PAD:18 PAD:32 0.586956
rPAD/11505 PAD:18 PAD:30 0.586956
rPAD/11506 PAD:18 PAD:9486 0.586956
rPAD/11507 PAD:18 PAD:9476 0.586956
rPAD/11508 PAD:18 PAD:9465 0.586956
rPAD/11509 PAD:18 PAD:9454 0.586956
rPAD/11510 PAD:18 PAD:19 0.9
rPAD/11511 R7:pos PAD:9423 0.0184795
rPAD/11512 R6:pos PAD:9410 0.0184795
rPAD/11513 R5:pos PAD:9397 0.0184795
rPAD/11514 R4:pos PAD:9387 0.0184795
rPAD/11515 R3:pos PAD:9370 0.0184795
rPAD/11516 R2:pos PAD:9358 0.0184795
rPAD/11517 R1:pos PAD:9345 0.0184795
rPAD/11518 R0:pos PAD:9332 0.0184795
cASIG5V/0 ASIG5V vss 73.974f
cASIG5V/1 ASIG5V vss 76.9788f
cASIG5V/2 ASIG5V vss 71.7842f
cASIG5V/3 ASIG5V vss 73.8848f
cASIG5V/4 ASIG5V vss 73.914f
cASIG5V/5 ASIG5V vss 71.7842f
cASIG5V/6 ASIG5V vss 74.11f
cASIG5V/7 ASIG5V vss 73.974f
cASIG5V/8 ASIG5V:1383 vss 28.7583f
cASIG5V/9 ASIG5V:1369 vss 36.9812f
cASIG5V/10 ASIG5V:1367 vss 28.7641f
cASIG5V/11 ASIG5V:1353 vss 36.8883f
cASIG5V/12 ASIG5V:1351 vss 28.7583f
cASIG5V/13 ASIG5V:1337 vss 36.0371f
cASIG5V/14 ASIG5V:1335 vss 28.7295f
cASIG5V/15 ASIG5V:1321 vss 36.7911f
cASIG5V/16 ASIG5V:1319 vss 28.7295f
cASIG5V/17 ASIG5V:1305 vss 36.7911f
cASIG5V/18 ASIG5V:1303 vss 28.7583f
cASIG5V/19 ASIG5V:1289 vss 36.0371f
cASIG5V/20 ASIG5V:1287 vss 28.7596f
cASIG5V/21 ASIG5V:1273 vss 36.8821f
cASIG5V/22 ASIG5V:1271 vss 28.7583f
cASIG5V/23 ASIG5V:1257 vss 36.9812f
cASIG5V/24 X46/X33/D0:pos vss 2.87453f
cASIG5V/25 ASIG5V:768 vss 7.64287f
cASIG5V/26 ASIG5V:663 vss 7.77059f
cASIG5V/27 X46/X31/D0:pos vss 2.88048f
cASIG5V/28 ASIG5V:558 vss 7.75131f
cASIG5V/29 X46/X30/D0:pos vss 2.93548f
cASIG5V/30 ASIG5V:453 vss 7.58192f
cASIG5V/31 X46/X29/D0:neg vss 4.13411f
cASIG5V/32 ASIG5V:416 vss 6.51082f
cASIG5V/33 X46/X28/D0:neg vss 4.18183f
cASIG5V/34 ASIG5V:311 vss 6.54488f
cASIG5V/35 X46/X27/D0:neg vss 2.97197f
cASIG5V/36 ASIG5V:138 vss 7.73761f
cASIG5V/37 X46/X26/D0:neg vss 2.99591f
cASIG5V/38 ASIG5V:33 vss 7.52148f
lASIG5V/39 ASIG5V:3083 R7:neg 4.67374p 
rASIG5V/40 ASIG5V:3083 ASIG5V:1383 0.361332
rASIG5V/41 ASIG5V:1384 ASIG5V:1383 0.225
lASIG5V/42 ASIG5V:3081 ASIG5V:1381 3.67204p 
rASIG5V/43 ASIG5V:3081 ASIG5V:1383 0.283889
rASIG5V/44 ASIG5V:1382 ASIG5V:1381 0.225
lASIG5V/45 ASIG5V:3079 ASIG5V:1379 3.67204p 
rASIG5V/46 ASIG5V:3079 ASIG5V:1381 0.283889
rASIG5V/47 ASIG5V:1380 ASIG5V:1379 0.225
lASIG5V/48 ASIG5V:3077 ASIG5V:1377 3.67204p 
rASIG5V/49 ASIG5V:3077 ASIG5V:1379 0.283889
rASIG5V/50 ASIG5V:1378 ASIG5V:1377 0.225
lASIG5V/51 ASIG5V:3075 ASIG5V:1375 8.35625p 
rASIG5V/52 ASIG5V:3075 ASIG5V:1377 0.64603
rASIG5V/53 ASIG5V:1376 ASIG5V:1375 0.225
lASIG5V/54 ASIG5V:3073 ASIG5V:1373 3.67204p 
rASIG5V/55 ASIG5V:3073 ASIG5V:1375 0.283889
rASIG5V/56 ASIG5V:1374 ASIG5V:1373 0.225
lASIG5V/57 ASIG5V:3071 ASIG5V:1371 3.67204p 
rASIG5V/58 ASIG5V:3071 ASIG5V:1373 0.283889
rASIG5V/59 ASIG5V:1372 ASIG5V:1371 0.225
lASIG5V/60 ASIG5V:3069 ASIG5V:1369 3.67204p 
rASIG5V/61 ASIG5V:3069 ASIG5V:1371 0.283889
lASIG5V/62 ASIG5V:3067 ASIG5V 96.4828p 
rASIG5V/63 ASIG5V:3067 ASIG5V:1369 9.27884
rASIG5V/64 ASIG5V:1370 ASIG5V:1369 0.225
lASIG5V/65 ASIG5V:3065 R6:neg 4.81274p 
rASIG5V/66 ASIG5V:3065 ASIG5V:1367 0.363399
rASIG5V/67 ASIG5V:1368 ASIG5V:1367 0.225
lASIG5V/68 ASIG5V:3063 ASIG5V:1365 3.78125p 
rASIG5V/69 ASIG5V:3063 ASIG5V:1367 0.285513
rASIG5V/70 ASIG5V:1366 ASIG5V:1365 0.225
lASIG5V/71 ASIG5V:3061 ASIG5V:1363 3.78125p 
rASIG5V/72 ASIG5V:3061 ASIG5V:1365 0.285513
rASIG5V/73 ASIG5V:1364 ASIG5V:1363 0.225
lASIG5V/74 ASIG5V:3059 ASIG5V:1361 3.78125p 
rASIG5V/75 ASIG5V:3059 ASIG5V:1363 0.285513
rASIG5V/76 ASIG5V:1362 ASIG5V:1361 0.225
lASIG5V/77 ASIG5V:3057 ASIG5V:1359 8.60476p 
rASIG5V/78 ASIG5V:3057 ASIG5V:1361 0.649726
rASIG5V/79 ASIG5V:1360 ASIG5V:1359 0.225
lASIG5V/80 ASIG5V:3055 ASIG5V:1357 3.78125p 
rASIG5V/81 ASIG5V:3055 ASIG5V:1359 0.285513
rASIG5V/82 ASIG5V:1358 ASIG5V:1357 0.225
lASIG5V/83 ASIG5V:3053 ASIG5V:1355 3.78125p 
rASIG5V/84 ASIG5V:3053 ASIG5V:1357 0.285513
rASIG5V/85 ASIG5V:1356 ASIG5V:1355 0.225
lASIG5V/86 ASIG5V:3051 ASIG5V:1353 3.78125p 
rASIG5V/87 ASIG5V:3051 ASIG5V:1355 0.285513
lASIG5V/88 ASIG5V:3049 ASIG5V 95.7151p 
rASIG5V/89 ASIG5V:3049 ASIG5V:1353 9.41378
rASIG5V/90 ASIG5V:1354 ASIG5V:1353 0.225
lASIG5V/91 ASIG5V:3047 R5:neg 6.07088p 
rASIG5V/92 ASIG5V:3047 ASIG5V:1351 0.369277
rASIG5V/93 ASIG5V:1352 ASIG5V:1351 0.225
lASIG5V/94 ASIG5V:3045 ASIG5V:1349 4.76974p 
rASIG5V/95 ASIG5V:3045 ASIG5V:1351 0.290132
rASIG5V/96 ASIG5V:1350 ASIG5V:1349 0.225
lASIG5V/97 ASIG5V:3043 ASIG5V:1347 4.76974p 
rASIG5V/98 ASIG5V:3043 ASIG5V:1349 0.290132
rASIG5V/99 ASIG5V:1348 ASIG5V:1347 0.225
lASIG5V/100 ASIG5V:3041 ASIG5V:1345 4.76974p 
rASIG5V/101 ASIG5V:3041 ASIG5V:1347 0.290132
rASIG5V/102 ASIG5V:1346 ASIG5V:1345 0.225
lASIG5V/103 ASIG5V:3039 ASIG5V:1343 10.8542p 
rASIG5V/104 ASIG5V:3039 ASIG5V:1345 0.660235
rASIG5V/105 ASIG5V:1344 ASIG5V:1343 0.225
lASIG5V/106 ASIG5V:3037 ASIG5V:1341 4.76974p 
rASIG5V/107 ASIG5V:3037 ASIG5V:1343 0.290132
rASIG5V/108 ASIG5V:1342 ASIG5V:1341 0.225
lASIG5V/109 ASIG5V:3035 ASIG5V:1339 4.76974p 
rASIG5V/110 ASIG5V:3035 ASIG5V:1341 0.290132
rASIG5V/111 ASIG5V:1340 ASIG5V:1339 0.225
lASIG5V/112 ASIG5V:3033 ASIG5V:1337 4.76974p 
rASIG5V/113 ASIG5V:3033 ASIG5V:1339 0.290132
lASIG5V/114 ASIG5V:3031 ASIG5V 111.72p 
rASIG5V/115 ASIG5V:3031 ASIG5V:1337 9.12149
rASIG5V/116 ASIG5V:1338 ASIG5V:1337 0.225
lASIG5V/117 ASIG5V:3029 R4:neg 4.85504p 
rASIG5V/118 ASIG5V:3029 ASIG5V:1335 0.384905
rASIG5V/119 ASIG5V:1336 ASIG5V:1335 0.225
lASIG5V/120 ASIG5V:3027 ASIG5V:1333 3.81448p 
rASIG5V/121 ASIG5V:3027 ASIG5V:1335 0.30241
rASIG5V/122 ASIG5V:1334 ASIG5V:1333 0.225
lASIG5V/123 ASIG5V:3025 ASIG5V:1331 3.81448p 
rASIG5V/124 ASIG5V:3025 ASIG5V:1333 0.30241
rASIG5V/125 ASIG5V:1332 ASIG5V:1331 0.225
lASIG5V/126 ASIG5V:3023 ASIG5V:1329 3.81448p 
rASIG5V/127 ASIG5V:3023 ASIG5V:1331 0.30241
rASIG5V/128 ASIG5V:1330 ASIG5V:1329 0.225
lASIG5V/129 ASIG5V:3021 ASIG5V:1327 8.68038p 
rASIG5V/130 ASIG5V:3021 ASIG5V:1329 0.688177
rASIG5V/131 ASIG5V:1328 ASIG5V:1327 0.225
lASIG5V/132 ASIG5V:3019 ASIG5V:1325 3.81448p 
rASIG5V/133 ASIG5V:3019 ASIG5V:1327 0.30241
rASIG5V/134 ASIG5V:1326 ASIG5V:1325 0.225
lASIG5V/135 ASIG5V:3017 ASIG5V:1323 3.81448p 
rASIG5V/136 ASIG5V:3017 ASIG5V:1325 0.30241
rASIG5V/137 ASIG5V:1324 ASIG5V:1323 0.225
lASIG5V/138 ASIG5V:3015 ASIG5V:1321 3.81448p 
rASIG5V/139 ASIG5V:3015 ASIG5V:1323 0.30241
lASIG5V/140 ASIG5V:3013 ASIG5V 111.621p 
rASIG5V/141 ASIG5V:3013 ASIG5V:1321 8.9712
rASIG5V/142 ASIG5V:1322 ASIG5V:1321 0.225
lASIG5V/143 ASIG5V:3011 R3:neg 4.9324p 
rASIG5V/144 ASIG5V:3011 ASIG5V:1319 0.38585
rASIG5V/145 ASIG5V:1320 ASIG5V:1319 0.225
lASIG5V/146 ASIG5V:3009 ASIG5V:1317 3.87526p 
rASIG5V/147 ASIG5V:3009 ASIG5V:1319 0.303152
rASIG5V/148 ASIG5V:1318 ASIG5V:1317 0.225
lASIG5V/149 ASIG5V:3007 ASIG5V:1315 3.87526p 
rASIG5V/150 ASIG5V:3007 ASIG5V:1317 0.303152
rASIG5V/151 ASIG5V:1316 ASIG5V:1315 0.225
lASIG5V/152 ASIG5V:3005 ASIG5V:1313 3.87526p 
rASIG5V/153 ASIG5V:3005 ASIG5V:1315 0.303152
rASIG5V/154 ASIG5V:1314 ASIG5V:1313 0.225
lASIG5V/155 ASIG5V:3003 ASIG5V:1311 8.8187p 
rASIG5V/156 ASIG5V:3003 ASIG5V:1313 0.689866
rASIG5V/157 ASIG5V:1312 ASIG5V:1311 0.225
lASIG5V/158 ASIG5V:3001 ASIG5V:1309 3.87526p 
rASIG5V/159 ASIG5V:3001 ASIG5V:1311 0.303152
rASIG5V/160 ASIG5V:1310 ASIG5V:1309 0.225
lASIG5V/161 ASIG5V:2999 ASIG5V:1307 3.87526p 
rASIG5V/162 ASIG5V:2999 ASIG5V:1309 0.303152
rASIG5V/163 ASIG5V:1308 ASIG5V:1307 0.225
lASIG5V/164 ASIG5V:2997 ASIG5V:1305 3.87526p 
rASIG5V/165 ASIG5V:2997 ASIG5V:1307 0.303152
lASIG5V/166 ASIG5V:2995 ASIG5V 118.329p 
rASIG5V/167 ASIG5V:2995 ASIG5V:1305 8.96285
rASIG5V/168 ASIG5V:1306 ASIG5V:1305 0.225
lASIG5V/169 ASIG5V:2993 R2:neg 4.86713p 
rASIG5V/170 ASIG5V:2993 ASIG5V:1303 0.364573
rASIG5V/171 ASIG5V:1304 ASIG5V:1303 0.225
lASIG5V/172 ASIG5V:2991 ASIG5V:1301 3.82398p 
rASIG5V/173 ASIG5V:2991 ASIG5V:1303 0.286436
rASIG5V/174 ASIG5V:1302 ASIG5V:1301 0.225
lASIG5V/175 ASIG5V:2989 ASIG5V:1299 3.82398p 
rASIG5V/176 ASIG5V:2989 ASIG5V:1301 0.286436
rASIG5V/177 ASIG5V:1300 ASIG5V:1299 0.225
lASIG5V/178 ASIG5V:2987 ASIG5V:1297 3.82398p 
rASIG5V/179 ASIG5V:2987 ASIG5V:1299 0.286436
rASIG5V/180 ASIG5V:1298 ASIG5V:1297 0.225
lASIG5V/181 ASIG5V:2985 ASIG5V:1295 8.70201p 
rASIG5V/182 ASIG5V:2985 ASIG5V:1297 0.651825
rASIG5V/183 ASIG5V:1296 ASIG5V:1295 0.225
lASIG5V/184 ASIG5V:2983 ASIG5V:1293 3.82398p 
rASIG5V/185 ASIG5V:2983 ASIG5V:1295 0.286436
rASIG5V/186 ASIG5V:1294 ASIG5V:1293 0.225
lASIG5V/187 ASIG5V:2981 ASIG5V:1291 3.82398p 
rASIG5V/188 ASIG5V:2981 ASIG5V:1293 0.286436
rASIG5V/189 ASIG5V:1292 ASIG5V:1291 0.225
lASIG5V/190 ASIG5V:2979 ASIG5V:1289 3.82398p 
rASIG5V/191 ASIG5V:2979 ASIG5V:1291 0.286436
lASIG5V/192 ASIG5V:2977 ASIG5V 118.347p 
rASIG5V/193 ASIG5V:2977 ASIG5V:1289 9.11067
rASIG5V/194 ASIG5V:1290 ASIG5V:1289 0.225
lASIG5V/195 ASIG5V:2975 R1:neg 4.5083p 
rASIG5V/196 ASIG5V:2975 ASIG5V:1287 0.362756
rASIG5V/197 ASIG5V:1288 ASIG5V:1287 0.225
lASIG5V/198 ASIG5V:2973 ASIG5V:1285 3.54206p 
rASIG5V/199 ASIG5V:2973 ASIG5V:1287 0.285008
rASIG5V/200 ASIG5V:1286 ASIG5V:1285 0.225
lASIG5V/201 ASIG5V:2971 ASIG5V:1283 3.54206p 
rASIG5V/202 ASIG5V:2971 ASIG5V:1285 0.285008
rASIG5V/203 ASIG5V:1284 ASIG5V:1283 0.225
lASIG5V/204 ASIG5V:2969 ASIG5V:1281 3.54206p 
rASIG5V/205 ASIG5V:2969 ASIG5V:1283 0.285008
rASIG5V/206 ASIG5V:1282 ASIG5V:1281 0.225
lASIG5V/207 ASIG5V:2967 ASIG5V:1279 8.06045p 
rASIG5V/208 ASIG5V:2967 ASIG5V:1281 0.648575
rASIG5V/209 ASIG5V:1280 ASIG5V:1279 0.225
lASIG5V/210 ASIG5V:2965 ASIG5V:1277 3.54206p 
rASIG5V/211 ASIG5V:2965 ASIG5V:1279 0.285008
rASIG5V/212 ASIG5V:1278 ASIG5V:1277 0.225
lASIG5V/213 ASIG5V:2963 ASIG5V:1275 3.54206p 
rASIG5V/214 ASIG5V:2963 ASIG5V:1277 0.285008
rASIG5V/215 ASIG5V:1276 ASIG5V:1275 0.225
lASIG5V/216 ASIG5V:2961 ASIG5V:1273 3.54206p 
rASIG5V/217 ASIG5V:2961 ASIG5V:1275 0.285008
lASIG5V/218 ASIG5V:2959 ASIG5V 102.413p 
rASIG5V/219 ASIG5V:2959 ASIG5V:1273 9.39452
rASIG5V/220 ASIG5V:1274 ASIG5V:1273 0.225
lASIG5V/221 ASIG5V:2957 R0:neg 4.38046p 
rASIG5V/222 ASIG5V:2957 ASIG5V:1271 0.361051
rASIG5V/223 ASIG5V:1272 ASIG5V:1271 0.225
lASIG5V/224 ASIG5V:2955 ASIG5V:1269 3.44162p 
rASIG5V/225 ASIG5V:2955 ASIG5V:1271 0.283668
rASIG5V/226 ASIG5V:1270 ASIG5V:1269 0.225
lASIG5V/227 ASIG5V:2953 ASIG5V:1267 3.44162p 
rASIG5V/228 ASIG5V:2953 ASIG5V:1269 0.283668
rASIG5V/229 ASIG5V:1268 ASIG5V:1267 0.225
lASIG5V/230 ASIG5V:2951 ASIG5V:1265 3.44162p 
rASIG5V/231 ASIG5V:2951 ASIG5V:1267 0.283668
rASIG5V/232 ASIG5V:1266 ASIG5V:1265 0.225
lASIG5V/233 ASIG5V:2949 ASIG5V:1263 7.83188p 
rASIG5V/234 ASIG5V:2949 ASIG5V:1265 0.645527
rASIG5V/235 ASIG5V:1264 ASIG5V:1263 0.225
lASIG5V/236 ASIG5V:2947 ASIG5V:1261 3.44162p 
rASIG5V/237 ASIG5V:2947 ASIG5V:1263 0.283668
rASIG5V/238 ASIG5V:1262 ASIG5V:1261 0.225
lASIG5V/239 ASIG5V:2945 ASIG5V:1259 3.44162p 
rASIG5V/240 ASIG5V:2945 ASIG5V:1261 0.283668
rASIG5V/241 ASIG5V:1260 ASIG5V:1259 0.225
lASIG5V/242 ASIG5V:2943 ASIG5V:1257 3.44162p 
rASIG5V/243 ASIG5V:2943 ASIG5V:1259 0.283668
lASIG5V/244 ASIG5V:2941 ASIG5V 99.8948p 
rASIG5V/245 ASIG5V:2941 ASIG5V:1257 9.21806
rASIG5V/246 ASIG5V:1258 ASIG5V:1257 0.225
rASIG5V/247 X46/X33/D0:pos ASIG5V:1378 0.445714
lASIG5V/248 ASIG5V:2939 ASIG5V:836 749.766f 
rASIG5V/249 ASIG5V:2939 ASIG5V:1378 0.0463984
rASIG5V/250 X46/X33/D0:pos ASIG5V:836 0.445714
rASIG5V/251 X46/X33/D0:pos ASIG5V:834 0.445714
lASIG5V/252 ASIG5V:2937 ASIG5V:832 514.303f 
rASIG5V/253 ASIG5V:2937 ASIG5V:1362 0.031827
rASIG5V/254 X46/X33/D0:pos ASIG5V:832 0.445714
rASIG5V/255 X46/X33/D0:pos ASIG5V:830 0.445714
lASIG5V/256 ASIG5V:2935 ASIG5V:828 285.035f 
rASIG5V/257 ASIG5V:2935 ASIG5V:1346 0.0176391
rASIG5V/258 X46/X33/D0:pos ASIG5V:828 0.445714
rASIG5V/259 X46/X33/D0:pos ASIG5V:826 0.445714
lASIG5V/260 ASIG5V:2933 ASIG5V:824 396.571f 
rASIG5V/261 ASIG5V:2933 ASIG5V:1330 0.0245413
rASIG5V/262 X46/X33/D0:pos ASIG5V:824 0.445714
rASIG5V/263 X46/X33/D0:pos ASIG5V:822 0.445714
rASIG5V/264 ASIG5V:820 X46/X33/D0:pos 0.445714
lASIG5V/265 ASIG5V:2931 ASIG5V:1314 408.963f 
rASIG5V/266 ASIG5V:2931 ASIG5V:818 0.0253082
rASIG5V/267 ASIG5V:818 X46/X33/D0:pos 0.445714
rASIG5V/268 ASIG5V:816 X46/X33/D0:pos 0.445714
lASIG5V/269 ASIG5V:2929 ASIG5V:1298 297.428f 
rASIG5V/270 ASIG5V:2929 ASIG5V:814 0.018406
rASIG5V/271 ASIG5V:814 X46/X33/D0:pos 0.445714
rASIG5V/272 ASIG5V:812 X46/X33/D0:pos 0.445714
lASIG5V/273 ASIG5V:2927 ASIG5V:1282 495.713f 
rASIG5V/274 ASIG5V:2927 ASIG5V:810 0.0306767
rASIG5V/275 ASIG5V:810 X46/X33/D0:pos 0.445714
rASIG5V/276 ASIG5V:808 X46/X33/D0:pos 0.445714
rASIG5V/277 ASIG5V:806 X46/X33/D0:pos 0.445714
lASIG5V/278 ASIG5V:2925 ASIG5V:834 625.838f 
rASIG5V/279 ASIG5V:2925 ASIG5V:800 0.0387293
rASIG5V/280 X46/X33/D0:pos ASIG5V:800 0.445714
lASIG5V/281 ASIG5V:2923 ASIG5V:1362 111.535f 
rASIG5V/282 ASIG5V:2923 ASIG5V:798 0.00690225
rASIG5V/283 X46/X33/D0:pos ASIG5V:798 0.445714
lASIG5V/284 ASIG5V:2921 ASIG5V:830 625.838f 
rASIG5V/285 ASIG5V:2921 ASIG5V:796 0.0387293
rASIG5V/286 X46/X33/D0:pos ASIG5V:796 0.445714
lASIG5V/287 ASIG5V:2919 ASIG5V:1346 24.7857f 
rASIG5V/288 ASIG5V:2919 ASIG5V:794 0.00153383
rASIG5V/289 X46/X33/D0:pos ASIG5V:794 0.445714
lASIG5V/290 ASIG5V:2917 ASIG5V:826 619.642f 
rASIG5V/291 ASIG5V:2917 ASIG5V:792 0.0383458
rASIG5V/292 X46/X33/D0:pos ASIG5V:792 0.445714
lASIG5V/293 ASIG5V:2915 ASIG5V:1330 223.071f 
rASIG5V/294 ASIG5V:2915 ASIG5V:790 0.0138045
rASIG5V/295 X46/X33/D0:pos ASIG5V:790 0.445714
lASIG5V/296 ASIG5V:2913 ASIG5V:822 619.642f 
rASIG5V/297 ASIG5V:2913 ASIG5V:788 0.0383458
rASIG5V/298 X46/X33/D0:pos ASIG5V:788 0.445714
lASIG5V/299 ASIG5V:2911 ASIG5V:820 619.642f 
rASIG5V/300 ASIG5V:2911 ASIG5V:786 0.0383458
rASIG5V/301 ASIG5V:786 X46/X33/D0:pos 0.445714
lASIG5V/302 ASIG5V:2909 ASIG5V:818 619.642f 
rASIG5V/303 ASIG5V:2909 ASIG5V:784 0.0383458
rASIG5V/304 ASIG5V:784 X46/X33/D0:pos 0.445714
lASIG5V/305 ASIG5V:2907 ASIG5V:816 309.821f 
rASIG5V/306 ASIG5V:2907 ASIG5V:782 0.0191729
rASIG5V/307 ASIG5V:782 X46/X33/D0:pos 0.445714
lASIG5V/308 ASIG5V:2905 ASIG5V:814 619.642f 
rASIG5V/309 ASIG5V:2905 ASIG5V:780 0.0383458
rASIG5V/310 ASIG5V:780 X46/X33/D0:pos 0.445714
lASIG5V/311 ASIG5V:2903 ASIG5V:812 619.642f 
rASIG5V/312 ASIG5V:2903 ASIG5V:778 0.0383458
rASIG5V/313 ASIG5V:778 X46/X33/D0:pos 0.445714
lASIG5V/314 ASIG5V:2901 ASIG5V:810 619.642f 
rASIG5V/315 ASIG5V:2901 ASIG5V:776 0.0383458
rASIG5V/316 ASIG5V:776 X46/X33/D0:pos 0.445714
lASIG5V/317 ASIG5V:2899 ASIG5V:774 545.285f 
rASIG5V/318 ASIG5V:2899 ASIG5V:1266 0.0337443
lASIG5V/319 ASIG5V:2897 ASIG5V:808 619.642f 
rASIG5V/320 ASIG5V:2897 ASIG5V:774 0.0383458
rASIG5V/321 ASIG5V:774 X46/X33/D0:pos 0.445714
lASIG5V/322 ASIG5V:2895 ASIG5V:806 619.642f 
rASIG5V/323 ASIG5V:2895 ASIG5V:772 0.0383458
rASIG5V/324 ASIG5V:772 X46/X33/D0:pos 0.445714
lASIG5V/325 ASIG5V:2893 X46/X33/D0:pos 619.642f 
rASIG5V/326 ASIG5V:2893 ASIG5V:772 0.352049
lASIG5V/327 ASIG5V:2891 ASIG5V:768 625.838f 
rASIG5V/328 ASIG5V:2891 ASIG5V:836 0.0387293
lASIG5V/329 ASIG5V:2889 ASIG5V:768 625.838f 
rASIG5V/330 ASIG5V:2889 X46/X33/D0:pos 0.270865
rASIG5V/331 X46/X33/D0:pos ASIG5V:768 0.445714
lASIG5V/332 ASIG5V:2887 ASIG5V:766 625.838f 
rASIG5V/333 ASIG5V:2887 ASIG5V:834 0.0387293
lASIG5V/334 ASIG5V:2885 ASIG5V:1378 501.91f 
rASIG5V/335 ASIG5V:2885 ASIG5V:766 0.0310601
rASIG5V/336 X46/X33/D0:pos ASIG5V:766 0.445714
lASIG5V/337 ASIG5V:2883 ASIG5V:764 625.838f 
rASIG5V/338 ASIG5V:2883 ASIG5V:832 0.0387293
lASIG5V/339 ASIG5V:2881 ASIG5V:800 625.838f 
rASIG5V/340 ASIG5V:2881 ASIG5V:764 0.0387293
rASIG5V/341 X46/X33/D0:pos ASIG5V:764 0.445714
lASIG5V/342 ASIG5V:2879 ASIG5V:762 625.838f 
rASIG5V/343 ASIG5V:2879 ASIG5V:830 0.0387293
lASIG5V/344 ASIG5V:2877 ASIG5V:798 625.838f 
rASIG5V/345 ASIG5V:2877 ASIG5V:762 0.0387293
rASIG5V/346 X46/X33/D0:pos ASIG5V:762 0.445714
lASIG5V/347 ASIG5V:2875 ASIG5V:760 619.642f 
rASIG5V/348 ASIG5V:2875 ASIG5V:828 0.0383458
lASIG5V/349 ASIG5V:2873 ASIG5V:796 625.838f 
rASIG5V/350 ASIG5V:2873 ASIG5V:760 0.0387293
rASIG5V/351 X46/X33/D0:pos ASIG5V:760 0.445714
lASIG5V/352 ASIG5V:2871 ASIG5V:758 309.821f 
rASIG5V/353 ASIG5V:2871 ASIG5V:826 0.0191729
lASIG5V/354 ASIG5V:2869 ASIG5V:794 929.462f 
rASIG5V/355 ASIG5V:2869 ASIG5V:758 0.0575187
rASIG5V/356 X46/X33/D0:pos ASIG5V:758 0.445714
lASIG5V/357 ASIG5V:2867 ASIG5V:756 619.642f 
rASIG5V/358 ASIG5V:2867 ASIG5V:824 0.0383458
lASIG5V/359 ASIG5V:2865 ASIG5V:792 619.642f 
rASIG5V/360 ASIG5V:2865 ASIG5V:756 0.0383458
rASIG5V/361 X46/X33/D0:pos ASIG5V:756 0.445714
lASIG5V/362 ASIG5V:2863 ASIG5V:754 619.642f 
rASIG5V/363 ASIG5V:2863 ASIG5V:822 0.0383458
lASIG5V/364 ASIG5V:2861 ASIG5V:790 619.642f 
rASIG5V/365 ASIG5V:2861 ASIG5V:754 0.0383458
rASIG5V/366 X46/X33/D0:pos ASIG5V:754 0.445714
lASIG5V/367 ASIG5V:2859 ASIG5V:752 619.642f 
rASIG5V/368 ASIG5V:2859 ASIG5V:820 0.0383458
lASIG5V/369 ASIG5V:2857 ASIG5V:788 619.642f 
rASIG5V/370 ASIG5V:2857 ASIG5V:752 0.0383458
rASIG5V/371 ASIG5V:752 X46/X33/D0:pos 0.445714
lASIG5V/372 ASIG5V:2855 ASIG5V:750 210.678f 
rASIG5V/373 ASIG5V:2855 ASIG5V:1314 0.0130376
lASIG5V/374 ASIG5V:2853 ASIG5V:786 619.642f 
rASIG5V/375 ASIG5V:2853 ASIG5V:750 0.0383458
rASIG5V/376 ASIG5V:750 X46/X33/D0:pos 0.445714
lASIG5V/377 ASIG5V:2851 ASIG5V:748 619.642f 
rASIG5V/378 ASIG5V:2851 ASIG5V:816 0.0383458
lASIG5V/379 ASIG5V:2849 ASIG5V:784 619.642f 
rASIG5V/380 ASIG5V:2849 ASIG5V:748 0.0383458
rASIG5V/381 ASIG5V:748 X46/X33/D0:pos 0.445714
lASIG5V/382 ASIG5V:2847 ASIG5V:746 12.3928f 
rASIG5V/383 ASIG5V:2847 ASIG5V:1298 0.000766916
lASIG5V/384 ASIG5V:2845 ASIG5V:782 929.462f 
rASIG5V/385 ASIG5V:2845 ASIG5V:746 0.0575187
rASIG5V/386 ASIG5V:746 X46/X33/D0:pos 0.445714
lASIG5V/387 ASIG5V:2843 ASIG5V:744 619.642f 
rASIG5V/388 ASIG5V:2843 ASIG5V:812 0.0383458
lASIG5V/389 ASIG5V:2841 ASIG5V:780 619.642f 
rASIG5V/390 ASIG5V:2841 ASIG5V:744 0.0383458
rASIG5V/391 ASIG5V:744 X46/X33/D0:pos 0.445714
lASIG5V/392 ASIG5V:2839 ASIG5V:742 123.928f 
rASIG5V/393 ASIG5V:2839 ASIG5V:1282 0.00766916
lASIG5V/394 ASIG5V:2837 ASIG5V:778 619.642f 
rASIG5V/395 ASIG5V:2837 ASIG5V:742 0.0383458
rASIG5V/396 ASIG5V:742 X46/X33/D0:pos 0.445714
lASIG5V/397 ASIG5V:2835 ASIG5V:740 619.642f 
rASIG5V/398 ASIG5V:2835 ASIG5V:808 0.0383458
lASIG5V/399 ASIG5V:2833 ASIG5V:776 619.642f 
rASIG5V/400 ASIG5V:2833 ASIG5V:740 0.0383458
rASIG5V/401 ASIG5V:740 X46/X33/D0:pos 0.445714
lASIG5V/402 ASIG5V:2831 ASIG5V:738 619.642f 
rASIG5V/403 ASIG5V:2831 ASIG5V:806 0.0383458
lASIG5V/404 ASIG5V:2829 ASIG5V:1266 74.357f 
rASIG5V/405 ASIG5V:2829 ASIG5V:738 0.0046015
rASIG5V/406 ASIG5V:738 X46/X33/D0:pos 0.445714
rASIG5V/407 X46/X32/D0:pos ASIG5V:1380 0.445714
lASIG5V/408 ASIG5V:2827 ASIG5V:731 856.274f 
rASIG5V/409 ASIG5V:2827 ASIG5V:1380 0.0444447
rASIG5V/410 X46/X32/D0:pos ASIG5V:731 0.445714
rASIG5V/411 X46/X32/D0:pos ASIG5V:729 0.445714
lASIG5V/412 ASIG5V:2825 ASIG5V:727 587.361f 
rASIG5V/413 ASIG5V:2825 ASIG5V:1364 0.0304869
rASIG5V/414 X46/X32/D0:pos ASIG5V:727 0.445714
rASIG5V/415 X46/X32/D0:pos ASIG5V:725 0.445714
lASIG5V/416 ASIG5V:2823 ASIG5V:723 325.526f 
rASIG5V/417 ASIG5V:2823 ASIG5V:1348 0.0168963
rASIG5V/418 X46/X32/D0:pos ASIG5V:723 0.445714
rASIG5V/419 X46/X32/D0:pos ASIG5V:721 0.445714
lASIG5V/420 ASIG5V:2821 ASIG5V:719 452.905f 
rASIG5V/421 ASIG5V:2821 ASIG5V:1332 0.0235079
rASIG5V/422 X46/X32/D0:pos ASIG5V:719 0.445714
rASIG5V/423 X46/X32/D0:pos ASIG5V:717 0.445714
rASIG5V/424 ASIG5V:715 X46/X32/D0:pos 0.445714
lASIG5V/425 ASIG5V:2819 ASIG5V:1316 467.059f 
rASIG5V/426 ASIG5V:2819 ASIG5V:713 0.0242426
rASIG5V/427 ASIG5V:713 X46/X32/D0:pos 0.445714
rASIG5V/428 ASIG5V:711 X46/X32/D0:pos 0.445714
lASIG5V/429 ASIG5V:2817 ASIG5V:1300 339.679f 
rASIG5V/430 ASIG5V:2817 ASIG5V:709 0.017631
rASIG5V/431 ASIG5V:709 X46/X32/D0:pos 0.445714
rASIG5V/432 ASIG5V:707 X46/X32/D0:pos 0.445714
lASIG5V/433 ASIG5V:2815 ASIG5V:1284 566.132f 
rASIG5V/434 ASIG5V:2815 ASIG5V:705 0.0293849
rASIG5V/435 ASIG5V:705 X46/X32/D0:pos 0.445714
rASIG5V/436 ASIG5V:703 X46/X32/D0:pos 0.445714
rASIG5V/437 ASIG5V:701 X46/X32/D0:pos 0.445714
lASIG5V/438 ASIG5V:2813 ASIG5V:729 714.741f 
rASIG5V/439 ASIG5V:2813 ASIG5V:695 0.0370985
rASIG5V/440 X46/X32/D0:pos ASIG5V:695 0.445714
lASIG5V/441 ASIG5V:2811 ASIG5V:1364 127.38f 
rASIG5V/442 ASIG5V:2811 ASIG5V:693 0.00661161
rASIG5V/443 X46/X32/D0:pos ASIG5V:693 0.445714
lASIG5V/444 ASIG5V:2809 ASIG5V:725 714.741f 
rASIG5V/445 ASIG5V:2809 ASIG5V:691 0.0370985
rASIG5V/446 X46/X32/D0:pos ASIG5V:691 0.445714
lASIG5V/447 ASIG5V:2807 ASIG5V:1348 28.3066f 
rASIG5V/448 ASIG5V:2807 ASIG5V:689 0.00146925
rASIG5V/449 X46/X32/D0:pos ASIG5V:689 0.445714
lASIG5V/450 ASIG5V:2805 ASIG5V:721 707.664f 
rASIG5V/451 ASIG5V:2805 ASIG5V:687 0.0367312
rASIG5V/452 X46/X32/D0:pos ASIG5V:687 0.445714
lASIG5V/453 ASIG5V:2803 ASIG5V:1332 254.759f 
rASIG5V/454 ASIG5V:2803 ASIG5V:685 0.0132232
rASIG5V/455 X46/X32/D0:pos ASIG5V:685 0.445714
lASIG5V/456 ASIG5V:2801 ASIG5V:717 707.664f 
rASIG5V/457 ASIG5V:2801 ASIG5V:683 0.0367312
rASIG5V/458 X46/X32/D0:pos ASIG5V:683 0.445714
lASIG5V/459 ASIG5V:2799 ASIG5V:715 707.664f 
rASIG5V/460 ASIG5V:2799 ASIG5V:681 0.0367312
rASIG5V/461 ASIG5V:681 X46/X32/D0:pos 0.445714
lASIG5V/462 ASIG5V:2797 ASIG5V:713 707.664f 
rASIG5V/463 ASIG5V:2797 ASIG5V:679 0.0367312
rASIG5V/464 ASIG5V:679 X46/X32/D0:pos 0.445714
lASIG5V/465 ASIG5V:2795 ASIG5V:711 353.832f 
rASIG5V/466 ASIG5V:2795 ASIG5V:677 0.0183656
rASIG5V/467 ASIG5V:677 X46/X32/D0:pos 0.445714
lASIG5V/468 ASIG5V:2793 ASIG5V:709 707.664f 
rASIG5V/469 ASIG5V:2793 ASIG5V:675 0.0367312
rASIG5V/470 ASIG5V:675 X46/X32/D0:pos 0.445714
lASIG5V/471 ASIG5V:2791 ASIG5V:707 707.664f 
rASIG5V/472 ASIG5V:2791 ASIG5V:673 0.0367312
rASIG5V/473 ASIG5V:673 X46/X32/D0:pos 0.445714
lASIG5V/474 ASIG5V:2789 ASIG5V:705 707.664f 
rASIG5V/475 ASIG5V:2789 ASIG5V:671 0.0367312
rASIG5V/476 ASIG5V:671 X46/X32/D0:pos 0.445714
lASIG5V/477 ASIG5V:2787 ASIG5V:669 622.745f 
rASIG5V/478 ASIG5V:2787 ASIG5V:1268 0.0323234
lASIG5V/479 ASIG5V:2785 ASIG5V:703 707.664f 
rASIG5V/480 ASIG5V:2785 ASIG5V:669 0.0367312
rASIG5V/481 ASIG5V:669 X46/X32/D0:pos 0.445714
lASIG5V/482 ASIG5V:2783 ASIG5V:701 707.664f 
rASIG5V/483 ASIG5V:2783 ASIG5V:667 0.0367312
rASIG5V/484 ASIG5V:667 X46/X32/D0:pos 0.445714
lASIG5V/485 ASIG5V:2781 X46/X32/D0:pos 707.664f 
rASIG5V/486 ASIG5V:2781 ASIG5V:667 0.350364
lASIG5V/487 ASIG5V:2779 ASIG5V:663 714.741f 
rASIG5V/488 ASIG5V:2779 ASIG5V:731 0.0370985
lASIG5V/489 ASIG5V:2777 ASIG5V:663 714.741f 
rASIG5V/490 ASIG5V:2777 X46/X32/D0:pos 0.26886
rASIG5V/491 X46/X32/D0:pos ASIG5V:663 0.445714
lASIG5V/492 ASIG5V:2775 ASIG5V:661 714.741f 
rASIG5V/493 ASIG5V:2775 ASIG5V:729 0.0370985
lASIG5V/494 ASIG5V:2773 ASIG5V:1380 573.208f 
rASIG5V/495 ASIG5V:2773 ASIG5V:661 0.0297522
rASIG5V/496 X46/X32/D0:pos ASIG5V:661 0.445714
lASIG5V/497 ASIG5V:2771 ASIG5V:659 714.741f 
rASIG5V/498 ASIG5V:2771 ASIG5V:727 0.0370985
lASIG5V/499 ASIG5V:2769 ASIG5V:695 714.741f 
rASIG5V/500 ASIG5V:2769 ASIG5V:659 0.0370985
rASIG5V/501 X46/X32/D0:pos ASIG5V:659 0.445714
lASIG5V/502 ASIG5V:2767 ASIG5V:657 714.741f 
rASIG5V/503 ASIG5V:2767 ASIG5V:725 0.0370985
lASIG5V/504 ASIG5V:2765 ASIG5V:693 714.741f 
rASIG5V/505 ASIG5V:2765 ASIG5V:657 0.0370985
rASIG5V/506 X46/X32/D0:pos ASIG5V:657 0.445714
lASIG5V/507 ASIG5V:2763 ASIG5V:655 707.664f 
rASIG5V/508 ASIG5V:2763 ASIG5V:723 0.0367312
lASIG5V/509 ASIG5V:2761 ASIG5V:691 714.741f 
rASIG5V/510 ASIG5V:2761 ASIG5V:655 0.0370985
rASIG5V/511 X46/X32/D0:pos ASIG5V:655 0.445714
lASIG5V/512 ASIG5V:2759 ASIG5V:653 353.832f 
rASIG5V/513 ASIG5V:2759 ASIG5V:721 0.0183656
lASIG5V/514 ASIG5V:2757 ASIG5V:689 1.0615p 
rASIG5V/515 ASIG5V:2757 ASIG5V:653 0.0550968
rASIG5V/516 X46/X32/D0:pos ASIG5V:653 0.445714
lASIG5V/517 ASIG5V:2755 ASIG5V:651 707.664f 
rASIG5V/518 ASIG5V:2755 ASIG5V:719 0.0367312
lASIG5V/519 ASIG5V:2753 ASIG5V:687 707.664f 
rASIG5V/520 ASIG5V:2753 ASIG5V:651 0.0367312
rASIG5V/521 X46/X32/D0:pos ASIG5V:651 0.445714
lASIG5V/522 ASIG5V:2751 ASIG5V:649 707.664f 
rASIG5V/523 ASIG5V:2751 ASIG5V:717 0.0367312
lASIG5V/524 ASIG5V:2749 ASIG5V:685 707.664f 
rASIG5V/525 ASIG5V:2749 ASIG5V:649 0.0367312
rASIG5V/526 X46/X32/D0:pos ASIG5V:649 0.445714
lASIG5V/527 ASIG5V:2747 ASIG5V:647 707.664f 
rASIG5V/528 ASIG5V:2747 ASIG5V:715 0.0367312
lASIG5V/529 ASIG5V:2745 ASIG5V:683 707.664f 
rASIG5V/530 ASIG5V:2745 ASIG5V:647 0.0367312
rASIG5V/531 ASIG5V:647 X46/X32/D0:pos 0.445714
lASIG5V/532 ASIG5V:2743 ASIG5V:645 240.606f 
rASIG5V/533 ASIG5V:2743 ASIG5V:1316 0.0124886
lASIG5V/534 ASIG5V:2741 ASIG5V:681 707.664f 
rASIG5V/535 ASIG5V:2741 ASIG5V:645 0.0367312
rASIG5V/536 ASIG5V:645 X46/X32/D0:pos 0.445714
lASIG5V/537 ASIG5V:2739 ASIG5V:643 707.664f 
rASIG5V/538 ASIG5V:2739 ASIG5V:711 0.0367312
lASIG5V/539 ASIG5V:2737 ASIG5V:679 707.664f 
rASIG5V/540 ASIG5V:2737 ASIG5V:643 0.0367312
rASIG5V/541 ASIG5V:643 X46/X32/D0:pos 0.445714
lASIG5V/542 ASIG5V:2735 ASIG5V:641 14.1533f 
rASIG5V/543 ASIG5V:2735 ASIG5V:1300 0.000734623
lASIG5V/544 ASIG5V:2733 ASIG5V:677 1.0615p 
rASIG5V/545 ASIG5V:2733 ASIG5V:641 0.0550968
rASIG5V/546 ASIG5V:641 X46/X32/D0:pos 0.445714
lASIG5V/547 ASIG5V:2731 ASIG5V:639 707.664f 
rASIG5V/548 ASIG5V:2731 ASIG5V:707 0.0367312
lASIG5V/549 ASIG5V:2729 ASIG5V:675 707.664f 
rASIG5V/550 ASIG5V:2729 ASIG5V:639 0.0367312
rASIG5V/551 ASIG5V:639 X46/X32/D0:pos 0.445714
lASIG5V/552 ASIG5V:2727 ASIG5V:637 141.533f 
rASIG5V/553 ASIG5V:2727 ASIG5V:1284 0.00734623
lASIG5V/554 ASIG5V:2725 ASIG5V:673 707.664f 
rASIG5V/555 ASIG5V:2725 ASIG5V:637 0.0367312
rASIG5V/556 ASIG5V:637 X46/X32/D0:pos 0.445714
lASIG5V/557 ASIG5V:2723 ASIG5V:635 707.664f 
rASIG5V/558 ASIG5V:2723 ASIG5V:703 0.0367312
lASIG5V/559 ASIG5V:2721 ASIG5V:671 707.664f 
rASIG5V/560 ASIG5V:2721 ASIG5V:635 0.0367312
rASIG5V/561 ASIG5V:635 X46/X32/D0:pos 0.445714
lASIG5V/562 ASIG5V:2719 ASIG5V:633 707.664f 
rASIG5V/563 ASIG5V:2719 ASIG5V:701 0.0367312
lASIG5V/564 ASIG5V:2717 ASIG5V:1268 84.9197f 
rASIG5V/565 ASIG5V:2717 ASIG5V:633 0.00440774
rASIG5V/566 ASIG5V:633 X46/X32/D0:pos 0.445714
rASIG5V/567 X46/X31/D0:pos ASIG5V:1382 0.445714
lASIG5V/568 ASIG5V:2715 ASIG5V:626 864.691f 
rASIG5V/569 ASIG5V:2715 ASIG5V:1382 0.0449716
rASIG5V/570 X46/X31/D0:pos ASIG5V:626 0.445714
rASIG5V/571 X46/X31/D0:pos ASIG5V:624 0.445714
lASIG5V/572 ASIG5V:2713 ASIG5V:622 593.135f 
rASIG5V/573 ASIG5V:2713 ASIG5V:1366 0.0308483
rASIG5V/574 X46/X31/D0:pos ASIG5V:622 0.445714
rASIG5V/575 X46/X31/D0:pos ASIG5V:620 0.445714
lASIG5V/576 ASIG5V:2711 ASIG5V:618 328.725f 
rASIG5V/577 ASIG5V:2711 ASIG5V:1350 0.0170967
rASIG5V/578 X46/X31/D0:pos ASIG5V:618 0.445714
rASIG5V/579 X46/X31/D0:pos ASIG5V:616 0.445714
lASIG5V/580 ASIG5V:2709 ASIG5V:614 457.357f 
rASIG5V/581 ASIG5V:2709 ASIG5V:1334 0.0237867
rASIG5V/582 X46/X31/D0:pos ASIG5V:614 0.445714
rASIG5V/583 X46/X31/D0:pos ASIG5V:612 0.445714
rASIG5V/584 ASIG5V:610 X46/X31/D0:pos 0.445714
lASIG5V/585 ASIG5V:2707 ASIG5V:1318 471.65f 
rASIG5V/586 ASIG5V:2707 ASIG5V:608 0.02453
rASIG5V/587 ASIG5V:608 X46/X31/D0:pos 0.445714
rASIG5V/588 ASIG5V:606 X46/X31/D0:pos 0.445714
lASIG5V/589 ASIG5V:2705 ASIG5V:1302 343.018f 
rASIG5V/590 ASIG5V:2705 ASIG5V:604 0.01784
rASIG5V/591 ASIG5V:604 X46/X31/D0:pos 0.445714
rASIG5V/592 ASIG5V:602 X46/X31/D0:pos 0.445714
lASIG5V/593 ASIG5V:2703 ASIG5V:1286 571.696f 
rASIG5V/594 ASIG5V:2703 ASIG5V:600 0.0297333
rASIG5V/595 ASIG5V:600 X46/X31/D0:pos 0.445714
rASIG5V/596 ASIG5V:598 X46/X31/D0:pos 0.445714
rASIG5V/597 ASIG5V:596 X46/X31/D0:pos 0.445714
lASIG5V/598 ASIG5V:2701 ASIG5V:624 721.767f 
rASIG5V/599 ASIG5V:2701 ASIG5V:590 0.0375383
rASIG5V/600 X46/X31/D0:pos ASIG5V:590 0.445714
lASIG5V/601 ASIG5V:2699 ASIG5V:1366 128.632f 
rASIG5V/602 ASIG5V:2699 ASIG5V:588 0.00669
rASIG5V/603 X46/X31/D0:pos ASIG5V:588 0.445714
lASIG5V/604 ASIG5V:2697 ASIG5V:620 721.767f 
rASIG5V/605 ASIG5V:2697 ASIG5V:586 0.0375383
rASIG5V/606 X46/X31/D0:pos ASIG5V:586 0.445714
lASIG5V/607 ASIG5V:2695 ASIG5V:1350 28.5848f 
rASIG5V/608 ASIG5V:2695 ASIG5V:584 0.00148667
rASIG5V/609 X46/X31/D0:pos ASIG5V:584 0.445714
lASIG5V/610 ASIG5V:2693 ASIG5V:616 714.62f 
rASIG5V/611 ASIG5V:2693 ASIG5V:582 0.0371666
rASIG5V/612 X46/X31/D0:pos ASIG5V:582 0.445714
lASIG5V/613 ASIG5V:2691 ASIG5V:1334 257.263f 
rASIG5V/614 ASIG5V:2691 ASIG5V:580 0.01338
rASIG5V/615 X46/X31/D0:pos ASIG5V:580 0.445714
lASIG5V/616 ASIG5V:2689 ASIG5V:612 714.62f 
rASIG5V/617 ASIG5V:2689 ASIG5V:578 0.0371666
rASIG5V/618 X46/X31/D0:pos ASIG5V:578 0.445714
lASIG5V/619 ASIG5V:2687 ASIG5V:610 714.62f 
rASIG5V/620 ASIG5V:2687 ASIG5V:576 0.0371666
rASIG5V/621 ASIG5V:576 X46/X31/D0:pos 0.445714
lASIG5V/622 ASIG5V:2685 ASIG5V:608 714.62f 
rASIG5V/623 ASIG5V:2685 ASIG5V:574 0.0371666
rASIG5V/624 ASIG5V:574 X46/X31/D0:pos 0.445714
lASIG5V/625 ASIG5V:2683 ASIG5V:606 357.31f 
rASIG5V/626 ASIG5V:2683 ASIG5V:572 0.0185833
rASIG5V/627 ASIG5V:572 X46/X31/D0:pos 0.445714
lASIG5V/628 ASIG5V:2681 ASIG5V:604 714.62f 
rASIG5V/629 ASIG5V:2681 ASIG5V:570 0.0371666
rASIG5V/630 ASIG5V:570 X46/X31/D0:pos 0.445714
lASIG5V/631 ASIG5V:2679 ASIG5V:602 714.62f 
rASIG5V/632 ASIG5V:2679 ASIG5V:568 0.0371666
rASIG5V/633 ASIG5V:568 X46/X31/D0:pos 0.445714
lASIG5V/634 ASIG5V:2677 ASIG5V:600 714.62f 
rASIG5V/635 ASIG5V:2677 ASIG5V:566 0.0371666
rASIG5V/636 ASIG5V:566 X46/X31/D0:pos 0.445714
lASIG5V/637 ASIG5V:2675 ASIG5V:564 628.866f 
rASIG5V/638 ASIG5V:2675 ASIG5V:1270 0.0327067
lASIG5V/639 ASIG5V:2673 ASIG5V:598 714.62f 
rASIG5V/640 ASIG5V:2673 ASIG5V:564 0.0371666
rASIG5V/641 ASIG5V:564 X46/X31/D0:pos 0.445714
lASIG5V/642 ASIG5V:2671 ASIG5V:596 714.62f 
rASIG5V/643 ASIG5V:2671 ASIG5V:562 0.0371666
rASIG5V/644 ASIG5V:562 X46/X31/D0:pos 0.445714
lASIG5V/645 ASIG5V:2669 X46/X31/D0:pos 714.62f 
rASIG5V/646 ASIG5V:2669 ASIG5V:562 0.350818
lASIG5V/647 ASIG5V:2667 ASIG5V:558 721.767f 
rASIG5V/648 ASIG5V:2667 ASIG5V:626 0.0375383
lASIG5V/649 ASIG5V:2665 ASIG5V:558 721.767f 
rASIG5V/650 ASIG5V:2665 X46/X31/D0:pos 0.269401
rASIG5V/651 X46/X31/D0:pos ASIG5V:558 0.445714
lASIG5V/652 ASIG5V:2663 ASIG5V:556 721.767f 
rASIG5V/653 ASIG5V:2663 ASIG5V:624 0.0375383
lASIG5V/654 ASIG5V:2661 ASIG5V:1382 578.843f 
rASIG5V/655 ASIG5V:2661 ASIG5V:556 0.030105
rASIG5V/656 X46/X31/D0:pos ASIG5V:556 0.445714
lASIG5V/657 ASIG5V:2659 ASIG5V:554 721.767f 
rASIG5V/658 ASIG5V:2659 ASIG5V:622 0.0375383
lASIG5V/659 ASIG5V:2657 ASIG5V:590 721.767f 
rASIG5V/660 ASIG5V:2657 ASIG5V:554 0.0375383
rASIG5V/661 X46/X31/D0:pos ASIG5V:554 0.445714
lASIG5V/662 ASIG5V:2655 ASIG5V:552 721.767f 
rASIG5V/663 ASIG5V:2655 ASIG5V:620 0.0375383
lASIG5V/664 ASIG5V:2653 ASIG5V:588 721.767f 
rASIG5V/665 ASIG5V:2653 ASIG5V:552 0.0375383
rASIG5V/666 X46/X31/D0:pos ASIG5V:552 0.445714
lASIG5V/667 ASIG5V:2651 ASIG5V:550 714.62f 
rASIG5V/668 ASIG5V:2651 ASIG5V:618 0.0371666
lASIG5V/669 ASIG5V:2649 ASIG5V:586 721.767f 
rASIG5V/670 ASIG5V:2649 ASIG5V:550 0.0375383
rASIG5V/671 X46/X31/D0:pos ASIG5V:550 0.445714
lASIG5V/672 ASIG5V:2647 ASIG5V:548 357.31f 
rASIG5V/673 ASIG5V:2647 ASIG5V:616 0.0185833
lASIG5V/674 ASIG5V:2645 ASIG5V:584 1.07193p 
rASIG5V/675 ASIG5V:2645 ASIG5V:548 0.05575
rASIG5V/676 X46/X31/D0:pos ASIG5V:548 0.445714
lASIG5V/677 ASIG5V:2643 ASIG5V:546 714.62f 
rASIG5V/678 ASIG5V:2643 ASIG5V:614 0.0371666
lASIG5V/679 ASIG5V:2641 ASIG5V:582 714.62f 
rASIG5V/680 ASIG5V:2641 ASIG5V:546 0.0371666
rASIG5V/681 X46/X31/D0:pos ASIG5V:546 0.445714
lASIG5V/682 ASIG5V:2639 ASIG5V:544 714.62f 
rASIG5V/683 ASIG5V:2639 ASIG5V:612 0.0371666
lASIG5V/684 ASIG5V:2637 ASIG5V:580 714.62f 
rASIG5V/685 ASIG5V:2637 ASIG5V:544 0.0371666
rASIG5V/686 X46/X31/D0:pos ASIG5V:544 0.445714
lASIG5V/687 ASIG5V:2635 ASIG5V:542 714.62f 
rASIG5V/688 ASIG5V:2635 ASIG5V:610 0.0371666
lASIG5V/689 ASIG5V:2633 ASIG5V:578 714.62f 
rASIG5V/690 ASIG5V:2633 ASIG5V:542 0.0371666
rASIG5V/691 ASIG5V:542 X46/X31/D0:pos 0.445714
lASIG5V/692 ASIG5V:2631 ASIG5V:540 242.971f 
rASIG5V/693 ASIG5V:2631 ASIG5V:1318 0.0126367
lASIG5V/694 ASIG5V:2629 ASIG5V:576 714.62f 
rASIG5V/695 ASIG5V:2629 ASIG5V:540 0.0371666
rASIG5V/696 ASIG5V:540 X46/X31/D0:pos 0.445714
lASIG5V/697 ASIG5V:2627 ASIG5V:538 714.62f 
rASIG5V/698 ASIG5V:2627 ASIG5V:606 0.0371666
lASIG5V/699 ASIG5V:2625 ASIG5V:574 714.62f 
rASIG5V/700 ASIG5V:2625 ASIG5V:538 0.0371666
rASIG5V/701 ASIG5V:538 X46/X31/D0:pos 0.445714
lASIG5V/702 ASIG5V:2623 ASIG5V:536 14.2924f 
rASIG5V/703 ASIG5V:2623 ASIG5V:1302 0.000743333
lASIG5V/704 ASIG5V:2621 ASIG5V:572 1.07193p 
rASIG5V/705 ASIG5V:2621 ASIG5V:536 0.05575
rASIG5V/706 ASIG5V:536 X46/X31/D0:pos 0.445714
lASIG5V/707 ASIG5V:2619 ASIG5V:534 714.62f 
rASIG5V/708 ASIG5V:2619 ASIG5V:602 0.0371666
lASIG5V/709 ASIG5V:2617 ASIG5V:570 714.62f 
rASIG5V/710 ASIG5V:2617 ASIG5V:534 0.0371666
rASIG5V/711 ASIG5V:534 X46/X31/D0:pos 0.445714
lASIG5V/712 ASIG5V:2615 ASIG5V:532 142.924f 
rASIG5V/713 ASIG5V:2615 ASIG5V:1286 0.00743333
lASIG5V/714 ASIG5V:2613 ASIG5V:568 714.62f 
rASIG5V/715 ASIG5V:2613 ASIG5V:532 0.0371666
rASIG5V/716 ASIG5V:532 X46/X31/D0:pos 0.445714
lASIG5V/717 ASIG5V:2611 ASIG5V:530 714.62f 
rASIG5V/718 ASIG5V:2611 ASIG5V:598 0.0371666
lASIG5V/719 ASIG5V:2609 ASIG5V:566 714.62f 
rASIG5V/720 ASIG5V:2609 ASIG5V:530 0.0371666
rASIG5V/721 ASIG5V:530 X46/X31/D0:pos 0.445714
lASIG5V/722 ASIG5V:2607 ASIG5V:528 714.62f 
rASIG5V/723 ASIG5V:2607 ASIG5V:596 0.0371666
lASIG5V/724 ASIG5V:2605 ASIG5V:1270 85.7545f 
rASIG5V/725 ASIG5V:2605 ASIG5V:528 0.00446
rASIG5V/726 ASIG5V:528 X46/X31/D0:pos 0.445714
rASIG5V/727 X46/X30/D0:pos ASIG5V:1384 0.445714
lASIG5V/728 ASIG5V:2603 ASIG5V:521 765.459f 
rASIG5V/729 ASIG5V:2603 ASIG5V:1384 0.048112
rASIG5V/730 X46/X30/D0:pos ASIG5V:521 0.445714
rASIG5V/731 X46/X30/D0:pos ASIG5V:519 0.445714
lASIG5V/732 ASIG5V:2601 ASIG5V:517 525.067f 
rASIG5V/733 ASIG5V:2601 ASIG5V:1368 0.0330024
rASIG5V/734 X46/X30/D0:pos ASIG5V:517 0.445714
rASIG5V/735 X46/X30/D0:pos ASIG5V:515 0.445714
lASIG5V/736 ASIG5V:2599 ASIG5V:513 291.001f 
rASIG5V/737 ASIG5V:2599 ASIG5V:1352 0.0182905
rASIG5V/738 X46/X30/D0:pos ASIG5V:513 0.445714
rASIG5V/739 X46/X30/D0:pos ASIG5V:511 0.445714
lASIG5V/740 ASIG5V:2597 ASIG5V:509 404.871f 
rASIG5V/741 ASIG5V:2597 ASIG5V:1336 0.0254477
rASIG5V/742 X46/X30/D0:pos ASIG5V:509 0.445714
rASIG5V/743 X46/X30/D0:pos ASIG5V:507 0.445714
rASIG5V/744 ASIG5V:505 X46/X30/D0:pos 0.445714
lASIG5V/745 ASIG5V:2595 ASIG5V:1320 417.523f 
rASIG5V/746 ASIG5V:2595 ASIG5V:503 0.0262429
rASIG5V/747 ASIG5V:503 X46/X30/D0:pos 0.445714
rASIG5V/748 ASIG5V:501 X46/X30/D0:pos 0.445714
lASIG5V/749 ASIG5V:2593 ASIG5V:1304 303.653f 
rASIG5V/750 ASIG5V:2593 ASIG5V:499 0.0190857
rASIG5V/751 ASIG5V:499 X46/X30/D0:pos 0.445714
rASIG5V/752 ASIG5V:497 X46/X30/D0:pos 0.445714
lASIG5V/753 ASIG5V:2591 ASIG5V:1288 506.089f 
rASIG5V/754 ASIG5V:2591 ASIG5V:495 0.0318096
rASIG5V/755 ASIG5V:495 X46/X30/D0:pos 0.445714
rASIG5V/756 ASIG5V:493 X46/X30/D0:pos 0.445714
rASIG5V/757 ASIG5V:491 X46/X30/D0:pos 0.445714
lASIG5V/758 ASIG5V:2589 ASIG5V:519 638.937f 
rASIG5V/759 ASIG5V:2589 ASIG5V:485 0.0401596
rASIG5V/760 X46/X30/D0:pos ASIG5V:485 0.445714
lASIG5V/761 ASIG5V:2587 ASIG5V:1368 113.87f 
rASIG5V/762 ASIG5V:2587 ASIG5V:483 0.00715715
rASIG5V/763 X46/X30/D0:pos ASIG5V:483 0.445714
lASIG5V/764 ASIG5V:2585 ASIG5V:515 638.937f 
rASIG5V/765 ASIG5V:2585 ASIG5V:481 0.0401596
rASIG5V/766 X46/X30/D0:pos ASIG5V:481 0.445714
lASIG5V/767 ASIG5V:2583 ASIG5V:1352 25.3044f 
rASIG5V/768 ASIG5V:2583 ASIG5V:479 0.00159048
rASIG5V/769 X46/X30/D0:pos ASIG5V:479 0.445714
lASIG5V/770 ASIG5V:2581 ASIG5V:511 632.611f 
rASIG5V/771 ASIG5V:2581 ASIG5V:477 0.039762
rASIG5V/772 X46/X30/D0:pos ASIG5V:477 0.445714
lASIG5V/773 ASIG5V:2579 ASIG5V:1336 227.74f 
rASIG5V/774 ASIG5V:2579 ASIG5V:475 0.0143143
rASIG5V/775 X46/X30/D0:pos ASIG5V:475 0.445714
lASIG5V/776 ASIG5V:2577 ASIG5V:507 632.611f 
rASIG5V/777 ASIG5V:2577 ASIG5V:473 0.039762
rASIG5V/778 X46/X30/D0:pos ASIG5V:473 0.445714
lASIG5V/779 ASIG5V:2575 ASIG5V:505 632.611f 
rASIG5V/780 ASIG5V:2575 ASIG5V:471 0.039762
rASIG5V/781 ASIG5V:471 X46/X30/D0:pos 0.445714
lASIG5V/782 ASIG5V:2573 ASIG5V:503 632.611f 
rASIG5V/783 ASIG5V:2573 ASIG5V:469 0.039762
rASIG5V/784 ASIG5V:469 X46/X30/D0:pos 0.445714
lASIG5V/785 ASIG5V:2571 ASIG5V:501 316.305f 
rASIG5V/786 ASIG5V:2571 ASIG5V:467 0.019881
rASIG5V/787 ASIG5V:467 X46/X30/D0:pos 0.445714
lASIG5V/788 ASIG5V:2569 ASIG5V:499 632.611f 
rASIG5V/789 ASIG5V:2569 ASIG5V:465 0.039762
rASIG5V/790 ASIG5V:465 X46/X30/D0:pos 0.445714
lASIG5V/791 ASIG5V:2567 ASIG5V:497 632.611f 
rASIG5V/792 ASIG5V:2567 ASIG5V:463 0.039762
rASIG5V/793 ASIG5V:463 X46/X30/D0:pos 0.445714
lASIG5V/794 ASIG5V:2565 ASIG5V:495 632.611f 
rASIG5V/795 ASIG5V:2565 ASIG5V:461 0.039762
rASIG5V/796 ASIG5V:461 X46/X30/D0:pos 0.445714
lASIG5V/797 ASIG5V:2563 ASIG5V:459 556.698f 
rASIG5V/798 ASIG5V:2563 ASIG5V:1272 0.0349905
lASIG5V/799 ASIG5V:2561 ASIG5V:493 632.611f 
rASIG5V/800 ASIG5V:2561 ASIG5V:459 0.039762
rASIG5V/801 ASIG5V:459 X46/X30/D0:pos 0.445714
lASIG5V/802 ASIG5V:2559 ASIG5V:491 632.611f 
rASIG5V/803 ASIG5V:2559 ASIG5V:457 0.039762
rASIG5V/804 ASIG5V:457 X46/X30/D0:pos 0.445714
lASIG5V/805 ASIG5V:2557 X46/X30/D0:pos 632.611f 
rASIG5V/806 ASIG5V:2557 ASIG5V:457 0.353527
lASIG5V/807 ASIG5V:2555 ASIG5V:453 638.937f 
rASIG5V/808 ASIG5V:2555 ASIG5V:521 0.0401596
lASIG5V/809 ASIG5V:2553 ASIG5V:453 638.937f 
rASIG5V/810 ASIG5V:2553 X46/X30/D0:pos 0.272624
rASIG5V/811 X46/X30/D0:pos ASIG5V:453 0.445714
lASIG5V/812 ASIG5V:2551 ASIG5V:451 638.937f 
rASIG5V/813 ASIG5V:2551 ASIG5V:519 0.0401596
lASIG5V/814 ASIG5V:2549 ASIG5V:1384 512.415f 
rASIG5V/815 ASIG5V:2549 ASIG5V:451 0.0322072
rASIG5V/816 X46/X30/D0:pos ASIG5V:451 0.445714
lASIG5V/817 ASIG5V:2547 ASIG5V:449 638.937f 
rASIG5V/818 ASIG5V:2547 ASIG5V:517 0.0401596
lASIG5V/819 ASIG5V:2545 ASIG5V:485 638.937f 
rASIG5V/820 ASIG5V:2545 ASIG5V:449 0.0401596
rASIG5V/821 X46/X30/D0:pos ASIG5V:449 0.445714
lASIG5V/822 ASIG5V:2543 ASIG5V:447 638.937f 
rASIG5V/823 ASIG5V:2543 ASIG5V:515 0.0401596
lASIG5V/824 ASIG5V:2541 ASIG5V:483 638.937f 
rASIG5V/825 ASIG5V:2541 ASIG5V:447 0.0401596
rASIG5V/826 X46/X30/D0:pos ASIG5V:447 0.445714
lASIG5V/827 ASIG5V:2539 ASIG5V:445 632.611f 
rASIG5V/828 ASIG5V:2539 ASIG5V:513 0.039762
lASIG5V/829 ASIG5V:2537 ASIG5V:481 638.937f 
rASIG5V/830 ASIG5V:2537 ASIG5V:445 0.0401596
rASIG5V/831 X46/X30/D0:pos ASIG5V:445 0.445714
lASIG5V/832 ASIG5V:2535 ASIG5V:443 316.305f 
rASIG5V/833 ASIG5V:2535 ASIG5V:511 0.019881
lASIG5V/834 ASIG5V:2533 ASIG5V:479 948.916f 
rASIG5V/835 ASIG5V:2533 ASIG5V:443 0.0596429
rASIG5V/836 X46/X30/D0:pos ASIG5V:443 0.445714
lASIG5V/837 ASIG5V:2531 ASIG5V:441 632.611f 
rASIG5V/838 ASIG5V:2531 ASIG5V:509 0.039762
lASIG5V/839 ASIG5V:2529 ASIG5V:477 632.611f 
rASIG5V/840 ASIG5V:2529 ASIG5V:441 0.039762
rASIG5V/841 X46/X30/D0:pos ASIG5V:441 0.445714
lASIG5V/842 ASIG5V:2527 ASIG5V:439 632.611f 
rASIG5V/843 ASIG5V:2527 ASIG5V:507 0.039762
lASIG5V/844 ASIG5V:2525 ASIG5V:475 632.611f 
rASIG5V/845 ASIG5V:2525 ASIG5V:439 0.039762
rASIG5V/846 X46/X30/D0:pos ASIG5V:439 0.445714
lASIG5V/847 ASIG5V:2523 ASIG5V:437 632.611f 
rASIG5V/848 ASIG5V:2523 ASIG5V:505 0.039762
lASIG5V/849 ASIG5V:2521 ASIG5V:473 632.611f 
rASIG5V/850 ASIG5V:2521 ASIG5V:437 0.039762
rASIG5V/851 ASIG5V:437 X46/X30/D0:pos 0.445714
lASIG5V/852 ASIG5V:2519 ASIG5V:435 215.088f 
rASIG5V/853 ASIG5V:2519 ASIG5V:1320 0.0135191
lASIG5V/854 ASIG5V:2517 ASIG5V:471 632.611f 
rASIG5V/855 ASIG5V:2517 ASIG5V:435 0.039762
rASIG5V/856 ASIG5V:435 X46/X30/D0:pos 0.445714
lASIG5V/857 ASIG5V:2515 ASIG5V:433 632.611f 
rASIG5V/858 ASIG5V:2515 ASIG5V:501 0.039762
lASIG5V/859 ASIG5V:2513 ASIG5V:469 632.611f 
rASIG5V/860 ASIG5V:2513 ASIG5V:433 0.039762
rASIG5V/861 ASIG5V:433 X46/X30/D0:pos 0.445714
lASIG5V/862 ASIG5V:2511 ASIG5V:431 12.6522f 
rASIG5V/863 ASIG5V:2511 ASIG5V:1304 0.000795239
lASIG5V/864 ASIG5V:2509 ASIG5V:467 948.916f 
rASIG5V/865 ASIG5V:2509 ASIG5V:431 0.0596429
rASIG5V/866 ASIG5V:431 X46/X30/D0:pos 0.445714
lASIG5V/867 ASIG5V:2507 ASIG5V:429 632.611f 
rASIG5V/868 ASIG5V:2507 ASIG5V:497 0.039762
lASIG5V/869 ASIG5V:2505 ASIG5V:465 632.611f 
rASIG5V/870 ASIG5V:2505 ASIG5V:429 0.039762
rASIG5V/871 ASIG5V:429 X46/X30/D0:pos 0.445714
lASIG5V/872 ASIG5V:2503 ASIG5V:427 126.522f 
rASIG5V/873 ASIG5V:2503 ASIG5V:1288 0.00795239
lASIG5V/874 ASIG5V:2501 ASIG5V:463 632.611f 
rASIG5V/875 ASIG5V:2501 ASIG5V:427 0.039762
rASIG5V/876 ASIG5V:427 X46/X30/D0:pos 0.445714
lASIG5V/877 ASIG5V:2499 ASIG5V:425 632.611f 
rASIG5V/878 ASIG5V:2499 ASIG5V:493 0.039762
lASIG5V/879 ASIG5V:2497 ASIG5V:461 632.611f 
rASIG5V/880 ASIG5V:2497 ASIG5V:425 0.039762
rASIG5V/881 ASIG5V:425 X46/X30/D0:pos 0.445714
lASIG5V/882 ASIG5V:2495 ASIG5V:423 632.611f 
rASIG5V/883 ASIG5V:2495 ASIG5V:491 0.039762
lASIG5V/884 ASIG5V:2493 ASIG5V:1272 75.9133f 
rASIG5V/885 ASIG5V:2493 ASIG5V:423 0.00477144
rASIG5V/886 ASIG5V:423 X46/X30/D0:pos 0.445714
rASIG5V/887 X46/X29/D0:neg ASIG5V:1370 0.445714
lASIG5V/888 ASIG5V:2491 ASIG5V:416 508.117f 
rASIG5V/889 ASIG5V:2491 ASIG5V:1370 0.04239
rASIG5V/890 X46/X29/D0:neg ASIG5V:416 0.445714
lASIG5V/891 ASIG5V:2489 ASIG5V:416 424.131f 
rASIG5V/892 ASIG5V:2489 X46/X29/D0:neg 0.20226
rASIG5V/893 X46/X29/D0:neg ASIG5V:414 0.445714
lASIG5V/894 ASIG5V:2487 ASIG5V:412 348.543f 
rASIG5V/895 ASIG5V:2487 ASIG5V:1354 0.0290774
rASIG5V/896 X46/X29/D0:neg ASIG5V:412 0.445714
rASIG5V/897 X46/X29/D0:neg ASIG5V:410 0.445714
lASIG5V/898 ASIG5V:2485 ASIG5V:408 193.169f 
rASIG5V/899 ASIG5V:2485 ASIG5V:1338 0.0161152
rASIG5V/900 X46/X29/D0:neg ASIG5V:408 0.445714
rASIG5V/901 X46/X29/D0:neg ASIG5V:406 0.445714
lASIG5V/902 ASIG5V:2483 ASIG5V:404 268.756f 
rASIG5V/903 ASIG5V:2483 ASIG5V:1322 0.0224212
rASIG5V/904 X46/X29/D0:neg ASIG5V:404 0.445714
rASIG5V/905 X46/X29/D0:neg ASIG5V:402 0.445714
rASIG5V/906 ASIG5V:400 X46/X29/D0:neg 0.445714
lASIG5V/907 ASIG5V:2481 ASIG5V:1306 277.155f 
rASIG5V/908 ASIG5V:2481 ASIG5V:398 0.0231218
rASIG5V/909 ASIG5V:398 X46/X29/D0:neg 0.445714
rASIG5V/910 ASIG5V:396 X46/X29/D0:neg 0.445714
lASIG5V/911 ASIG5V:2479 ASIG5V:1290 201.567f 
rASIG5V/912 ASIG5V:2479 ASIG5V:394 0.0168159
rASIG5V/913 ASIG5V:394 X46/X29/D0:neg 0.445714
rASIG5V/914 ASIG5V:392 X46/X29/D0:neg 0.445714
lASIG5V/915 ASIG5V:2477 ASIG5V:1274 335.945f 
rASIG5V/916 ASIG5V:2477 ASIG5V:390 0.0280264
rASIG5V/917 ASIG5V:390 X46/X29/D0:neg 0.445714
rASIG5V/918 ASIG5V:388 X46/X29/D0:neg 0.445714
rASIG5V/919 ASIG5V:386 X46/X29/D0:neg 0.445714
lASIG5V/920 ASIG5V:2475 X46/X29/D0:neg 419.932f 
rASIG5V/921 ASIG5V:2475 ASIG5V:386 0.23064
lASIG5V/922 ASIG5V:2473 ASIG5V:414 424.131f 
rASIG5V/923 ASIG5V:2473 ASIG5V:380 0.0353834
rASIG5V/924 X46/X29/D0:neg ASIG5V:380 0.445714
lASIG5V/925 ASIG5V:2471 ASIG5V:1354 75.5877f 
rASIG5V/926 ASIG5V:2471 ASIG5V:378 0.00630595
rASIG5V/927 X46/X29/D0:neg ASIG5V:378 0.445714
lASIG5V/928 ASIG5V:2469 ASIG5V:410 424.131f 
rASIG5V/929 ASIG5V:2469 ASIG5V:376 0.0353834
rASIG5V/930 X46/X29/D0:neg ASIG5V:376 0.445714
lASIG5V/931 ASIG5V:2467 ASIG5V:1338 16.7973f 
rASIG5V/932 ASIG5V:2467 ASIG5V:374 0.00140132
rASIG5V/933 X46/X29/D0:neg ASIG5V:374 0.445714
lASIG5V/934 ASIG5V:2465 ASIG5V:406 419.932f 
rASIG5V/935 ASIG5V:2465 ASIG5V:372 0.0350331
rASIG5V/936 X46/X29/D0:neg ASIG5V:372 0.445714
lASIG5V/937 ASIG5V:2463 ASIG5V:1322 151.175f 
rASIG5V/938 ASIG5V:2463 ASIG5V:370 0.0126119
rASIG5V/939 X46/X29/D0:neg ASIG5V:370 0.445714
lASIG5V/940 ASIG5V:2461 ASIG5V:402 419.932f 
rASIG5V/941 ASIG5V:2461 ASIG5V:368 0.0350331
rASIG5V/942 X46/X29/D0:neg ASIG5V:368 0.445714
lASIG5V/943 ASIG5V:2459 ASIG5V:400 419.932f 
rASIG5V/944 ASIG5V:2459 ASIG5V:366 0.0350331
rASIG5V/945 ASIG5V:366 X46/X29/D0:neg 0.445714
lASIG5V/946 ASIG5V:2457 ASIG5V:398 419.932f 
rASIG5V/947 ASIG5V:2457 ASIG5V:364 0.0350331
rASIG5V/948 ASIG5V:364 X46/X29/D0:neg 0.445714
lASIG5V/949 ASIG5V:2455 ASIG5V:396 209.966f 
rASIG5V/950 ASIG5V:2455 ASIG5V:362 0.0175165
rASIG5V/951 ASIG5V:362 X46/X29/D0:neg 0.445714
lASIG5V/952 ASIG5V:2453 ASIG5V:394 419.932f 
rASIG5V/953 ASIG5V:2453 ASIG5V:360 0.0350331
rASIG5V/954 ASIG5V:360 X46/X29/D0:neg 0.445714
lASIG5V/955 ASIG5V:2451 ASIG5V:392 419.932f 
rASIG5V/956 ASIG5V:2451 ASIG5V:358 0.0350331
rASIG5V/957 ASIG5V:358 X46/X29/D0:neg 0.445714
lASIG5V/958 ASIG5V:2449 ASIG5V:390 419.932f 
rASIG5V/959 ASIG5V:2449 ASIG5V:356 0.0350331
rASIG5V/960 ASIG5V:356 X46/X29/D0:neg 0.445714
lASIG5V/961 ASIG5V:2447 ASIG5V:354 369.54f 
rASIG5V/962 ASIG5V:2447 ASIG5V:1258 0.0308291
lASIG5V/963 ASIG5V:2445 ASIG5V:388 419.932f 
rASIG5V/964 ASIG5V:2445 ASIG5V:354 0.0350331
rASIG5V/965 ASIG5V:354 X46/X29/D0:neg 0.445714
lASIG5V/966 ASIG5V:2443 ASIG5V:346 424.131f 
rASIG5V/967 ASIG5V:2443 ASIG5V:414 0.0353834
lASIG5V/968 ASIG5V:2441 ASIG5V:1370 340.145f 
rASIG5V/969 ASIG5V:2441 ASIG5V:346 0.0283768
rASIG5V/970 X46/X29/D0:neg ASIG5V:346 0.445714
lASIG5V/971 ASIG5V:2439 ASIG5V:344 424.131f 
rASIG5V/972 ASIG5V:2439 ASIG5V:412 0.0353834
lASIG5V/973 ASIG5V:2437 ASIG5V:380 424.131f 
rASIG5V/974 ASIG5V:2437 ASIG5V:344 0.0353834
rASIG5V/975 X46/X29/D0:neg ASIG5V:344 0.445714
lASIG5V/976 ASIG5V:2435 ASIG5V:342 424.131f 
rASIG5V/977 ASIG5V:2435 ASIG5V:410 0.0353834
lASIG5V/978 ASIG5V:2433 ASIG5V:378 424.131f 
rASIG5V/979 ASIG5V:2433 ASIG5V:342 0.0353834
rASIG5V/980 X46/X29/D0:neg ASIG5V:342 0.445714
lASIG5V/981 ASIG5V:2431 ASIG5V:340 419.932f 
rASIG5V/982 ASIG5V:2431 ASIG5V:408 0.0350331
lASIG5V/983 ASIG5V:2429 ASIG5V:376 424.131f 
rASIG5V/984 ASIG5V:2429 ASIG5V:340 0.0353834
rASIG5V/985 X46/X29/D0:neg ASIG5V:340 0.445714
lASIG5V/986 ASIG5V:2427 ASIG5V:338 209.966f 
rASIG5V/987 ASIG5V:2427 ASIG5V:406 0.0175165
lASIG5V/988 ASIG5V:2425 ASIG5V:374 629.898f 
rASIG5V/989 ASIG5V:2425 ASIG5V:338 0.0525496
rASIG5V/990 X46/X29/D0:neg ASIG5V:338 0.445714
lASIG5V/991 ASIG5V:2423 ASIG5V:336 419.932f 
rASIG5V/992 ASIG5V:2423 ASIG5V:404 0.0350331
lASIG5V/993 ASIG5V:2421 ASIG5V:372 419.932f 
rASIG5V/994 ASIG5V:2421 ASIG5V:336 0.0350331
rASIG5V/995 X46/X29/D0:neg ASIG5V:336 0.445714
lASIG5V/996 ASIG5V:2419 ASIG5V:334 419.932f 
rASIG5V/997 ASIG5V:2419 ASIG5V:402 0.0350331
lASIG5V/998 ASIG5V:2417 ASIG5V:370 419.932f 
rASIG5V/999 ASIG5V:2417 ASIG5V:334 0.0350331
rASIG5V/1000 X46/X29/D0:neg ASIG5V:334 0.445714
lASIG5V/1001 ASIG5V:2415 ASIG5V:332 419.932f 
rASIG5V/1002 ASIG5V:2415 ASIG5V:400 0.0350331
lASIG5V/1003 ASIG5V:2413 ASIG5V:368 419.932f 
rASIG5V/1004 ASIG5V:2413 ASIG5V:332 0.0350331
rASIG5V/1005 ASIG5V:332 X46/X29/D0:neg 0.445714
lASIG5V/1006 ASIG5V:2411 ASIG5V:330 142.777f 
rASIG5V/1007 ASIG5V:2411 ASIG5V:1306 0.0119112
lASIG5V/1008 ASIG5V:2409 ASIG5V:366 419.932f 
rASIG5V/1009 ASIG5V:2409 ASIG5V:330 0.0350331
rASIG5V/1010 ASIG5V:330 X46/X29/D0:neg 0.445714
lASIG5V/1011 ASIG5V:2407 ASIG5V:328 419.932f 
rASIG5V/1012 ASIG5V:2407 ASIG5V:396 0.0350331
lASIG5V/1013 ASIG5V:2405 ASIG5V:364 419.932f 
rASIG5V/1014 ASIG5V:2405 ASIG5V:328 0.0350331
rASIG5V/1015 ASIG5V:328 X46/X29/D0:neg 0.445714
lASIG5V/1016 ASIG5V:2403 ASIG5V:326 8.39864f 
rASIG5V/1017 ASIG5V:2403 ASIG5V:1290 0.000700661
lASIG5V/1018 ASIG5V:2401 ASIG5V:362 629.898f 
rASIG5V/1019 ASIG5V:2401 ASIG5V:326 0.0525496
rASIG5V/1020 ASIG5V:326 X46/X29/D0:neg 0.445714
lASIG5V/1021 ASIG5V:2399 ASIG5V:324 419.932f 
rASIG5V/1022 ASIG5V:2399 ASIG5V:392 0.0350331
lASIG5V/1023 ASIG5V:2397 ASIG5V:360 419.932f 
rASIG5V/1024 ASIG5V:2397 ASIG5V:324 0.0350331
rASIG5V/1025 ASIG5V:324 X46/X29/D0:neg 0.445714
lASIG5V/1026 ASIG5V:2395 ASIG5V:322 83.9864f 
rASIG5V/1027 ASIG5V:2395 ASIG5V:1274 0.00700661
lASIG5V/1028 ASIG5V:2393 ASIG5V:358 419.932f 
rASIG5V/1029 ASIG5V:2393 ASIG5V:322 0.0350331
rASIG5V/1030 ASIG5V:322 X46/X29/D0:neg 0.445714
lASIG5V/1031 ASIG5V:2391 ASIG5V:320 419.932f 
rASIG5V/1032 ASIG5V:2391 ASIG5V:388 0.0350331
lASIG5V/1033 ASIG5V:2389 ASIG5V:356 419.932f 
rASIG5V/1034 ASIG5V:2389 ASIG5V:320 0.0350331
rASIG5V/1035 ASIG5V:320 X46/X29/D0:neg 0.445714
lASIG5V/1036 ASIG5V:2387 ASIG5V:318 419.932f 
rASIG5V/1037 ASIG5V:2387 ASIG5V:386 0.0350331
lASIG5V/1038 ASIG5V:2385 ASIG5V:1258 50.3918f 
rASIG5V/1039 ASIG5V:2385 ASIG5V:318 0.00420397
rASIG5V/1040 ASIG5V:318 X46/X29/D0:neg 0.445714
rASIG5V/1041 X46/X28/D0:neg ASIG5V:1372 0.445714
lASIG5V/1042 ASIG5V:2383 ASIG5V:311 487.532f 
rASIG5V/1043 ASIG5V:2383 ASIG5V:1372 0.0422446
rASIG5V/1044 X46/X28/D0:neg ASIG5V:311 0.445714
lASIG5V/1045 ASIG5V:2381 ASIG5V:311 406.948f 
rASIG5V/1046 ASIG5V:2381 X46/X28/D0:neg 0.20208
rASIG5V/1047 X46/X28/D0:neg ASIG5V:309 0.445714
lASIG5V/1048 ASIG5V:2379 ASIG5V:307 334.423f 
rASIG5V/1049 ASIG5V:2379 ASIG5V:1356 0.0289777
rASIG5V/1050 X46/X28/D0:neg ASIG5V:307 0.445714
rASIG5V/1051 X46/X28/D0:neg ASIG5V:305 0.445714
lASIG5V/1052 ASIG5V:2377 ASIG5V:303 185.343f 
rASIG5V/1053 ASIG5V:2377 ASIG5V:1340 0.0160599
rASIG5V/1054 X46/X28/D0:neg ASIG5V:303 0.445714
rASIG5V/1055 X46/X28/D0:neg ASIG5V:301 0.445714
lASIG5V/1056 ASIG5V:2375 ASIG5V:299 257.868f 
rASIG5V/1057 ASIG5V:2375 ASIG5V:1324 0.0223443
rASIG5V/1058 X46/X28/D0:neg ASIG5V:299 0.445714
rASIG5V/1059 X46/X28/D0:neg ASIG5V:297 0.445714
rASIG5V/1060 ASIG5V:295 X46/X28/D0:neg 0.445714
lASIG5V/1061 ASIG5V:2373 ASIG5V:1308 265.926f 
rASIG5V/1062 ASIG5V:2373 ASIG5V:293 0.0230425
rASIG5V/1063 ASIG5V:293 X46/X28/D0:neg 0.445714
rASIG5V/1064 ASIG5V:291 X46/X28/D0:neg 0.445714
lASIG5V/1065 ASIG5V:2371 ASIG5V:1292 193.401f 
rASIG5V/1066 ASIG5V:2371 ASIG5V:289 0.0167582
rASIG5V/1067 ASIG5V:289 X46/X28/D0:neg 0.445714
rASIG5V/1068 ASIG5V:287 X46/X28/D0:neg 0.445714
lASIG5V/1069 ASIG5V:2369 ASIG5V:1276 322.335f 
rASIG5V/1070 ASIG5V:2369 ASIG5V:285 0.0279303
rASIG5V/1071 ASIG5V:285 X46/X28/D0:neg 0.445714
rASIG5V/1072 ASIG5V:283 X46/X28/D0:neg 0.445714
rASIG5V/1073 ASIG5V:281 X46/X28/D0:neg 0.445714
lASIG5V/1074 ASIG5V:2367 X46/X28/D0:neg 402.919f 
rASIG5V/1075 ASIG5V:2367 ASIG5V:281 0.230481
lASIG5V/1076 ASIG5V:2365 ASIG5V:309 406.948f 
rASIG5V/1077 ASIG5V:2365 ASIG5V:275 0.035262
rASIG5V/1078 X46/X28/D0:neg ASIG5V:275 0.445714
lASIG5V/1079 ASIG5V:2363 ASIG5V:1356 72.5254f 
rASIG5V/1080 ASIG5V:2363 ASIG5V:273 0.00628432
rASIG5V/1081 X46/X28/D0:neg ASIG5V:273 0.445714
lASIG5V/1082 ASIG5V:2361 ASIG5V:305 406.948f 
rASIG5V/1083 ASIG5V:2361 ASIG5V:271 0.035262
rASIG5V/1084 X46/X28/D0:neg ASIG5V:271 0.445714
lASIG5V/1085 ASIG5V:2359 ASIG5V:1340 16.1167f 
rASIG5V/1086 ASIG5V:2359 ASIG5V:269 0.00139652
rASIG5V/1087 X46/X28/D0:neg ASIG5V:269 0.445714
lASIG5V/1088 ASIG5V:2357 ASIG5V:301 402.919f 
rASIG5V/1089 ASIG5V:2357 ASIG5V:267 0.0349129
rASIG5V/1090 X46/X28/D0:neg ASIG5V:267 0.445714
lASIG5V/1091 ASIG5V:2355 ASIG5V:1324 145.051f 
rASIG5V/1092 ASIG5V:2355 ASIG5V:265 0.0125686
rASIG5V/1093 X46/X28/D0:neg ASIG5V:265 0.445714
lASIG5V/1094 ASIG5V:2353 ASIG5V:297 402.919f 
rASIG5V/1095 ASIG5V:2353 ASIG5V:263 0.0349129
rASIG5V/1096 X46/X28/D0:neg ASIG5V:263 0.445714
lASIG5V/1097 ASIG5V:2351 ASIG5V:295 402.919f 
rASIG5V/1098 ASIG5V:2351 ASIG5V:261 0.0349129
rASIG5V/1099 ASIG5V:261 X46/X28/D0:neg 0.445714
lASIG5V/1100 ASIG5V:2349 ASIG5V:293 402.919f 
rASIG5V/1101 ASIG5V:2349 ASIG5V:259 0.0349129
rASIG5V/1102 ASIG5V:259 X46/X28/D0:neg 0.445714
lASIG5V/1103 ASIG5V:2347 ASIG5V:291 201.459f 
rASIG5V/1104 ASIG5V:2347 ASIG5V:257 0.0174565
rASIG5V/1105 ASIG5V:257 X46/X28/D0:neg 0.445714
lASIG5V/1106 ASIG5V:2345 ASIG5V:289 402.919f 
rASIG5V/1107 ASIG5V:2345 ASIG5V:255 0.0349129
rASIG5V/1108 ASIG5V:255 X46/X28/D0:neg 0.445714
lASIG5V/1109 ASIG5V:2343 ASIG5V:287 402.919f 
rASIG5V/1110 ASIG5V:2343 ASIG5V:253 0.0349129
rASIG5V/1111 ASIG5V:253 X46/X28/D0:neg 0.445714
lASIG5V/1112 ASIG5V:2341 ASIG5V:285 402.919f 
rASIG5V/1113 ASIG5V:2341 ASIG5V:251 0.0349129
rASIG5V/1114 ASIG5V:251 X46/X28/D0:neg 0.445714
lASIG5V/1115 ASIG5V:2339 ASIG5V:249 354.568f 
rASIG5V/1116 ASIG5V:2339 ASIG5V:1260 0.0307234
lASIG5V/1117 ASIG5V:2337 ASIG5V:283 402.919f 
rASIG5V/1118 ASIG5V:2337 ASIG5V:249 0.0349129
rASIG5V/1119 ASIG5V:249 X46/X28/D0:neg 0.445714
lASIG5V/1120 ASIG5V:2335 ASIG5V:241 406.948f 
rASIG5V/1121 ASIG5V:2335 ASIG5V:309 0.035262
lASIG5V/1122 ASIG5V:2333 ASIG5V:1372 326.364f 
rASIG5V/1123 ASIG5V:2333 ASIG5V:241 0.0282795
rASIG5V/1124 X46/X28/D0:neg ASIG5V:241 0.445714
lASIG5V/1125 ASIG5V:2331 ASIG5V:239 406.948f 
rASIG5V/1126 ASIG5V:2331 ASIG5V:307 0.035262
lASIG5V/1127 ASIG5V:2329 ASIG5V:275 406.948f 
rASIG5V/1128 ASIG5V:2329 ASIG5V:239 0.035262
rASIG5V/1129 X46/X28/D0:neg ASIG5V:239 0.445714
lASIG5V/1130 ASIG5V:2327 ASIG5V:237 406.948f 
rASIG5V/1131 ASIG5V:2327 ASIG5V:305 0.035262
lASIG5V/1132 ASIG5V:2325 ASIG5V:273 406.948f 
rASIG5V/1133 ASIG5V:2325 ASIG5V:237 0.035262
rASIG5V/1134 X46/X28/D0:neg ASIG5V:237 0.445714
lASIG5V/1135 ASIG5V:2323 ASIG5V:235 402.919f 
rASIG5V/1136 ASIG5V:2323 ASIG5V:303 0.0349129
lASIG5V/1137 ASIG5V:2321 ASIG5V:271 406.948f 
rASIG5V/1138 ASIG5V:2321 ASIG5V:235 0.035262
rASIG5V/1139 X46/X28/D0:neg ASIG5V:235 0.445714
lASIG5V/1140 ASIG5V:2319 ASIG5V:233 201.459f 
rASIG5V/1141 ASIG5V:2319 ASIG5V:301 0.0174565
lASIG5V/1142 ASIG5V:2317 ASIG5V:269 604.378f 
rASIG5V/1143 ASIG5V:2317 ASIG5V:233 0.0523694
rASIG5V/1144 X46/X28/D0:neg ASIG5V:233 0.445714
lASIG5V/1145 ASIG5V:2315 ASIG5V:231 402.919f 
rASIG5V/1146 ASIG5V:2315 ASIG5V:299 0.0349129
lASIG5V/1147 ASIG5V:2313 ASIG5V:267 402.919f 
rASIG5V/1148 ASIG5V:2313 ASIG5V:231 0.0349129
rASIG5V/1149 X46/X28/D0:neg ASIG5V:231 0.445714
lASIG5V/1150 ASIG5V:2311 ASIG5V:229 402.919f 
rASIG5V/1151 ASIG5V:2311 ASIG5V:297 0.0349129
lASIG5V/1152 ASIG5V:2309 ASIG5V:265 402.919f 
rASIG5V/1153 ASIG5V:2309 ASIG5V:229 0.0349129
rASIG5V/1154 X46/X28/D0:neg ASIG5V:229 0.445714
lASIG5V/1155 ASIG5V:2307 ASIG5V:227 402.919f 
rASIG5V/1156 ASIG5V:2307 ASIG5V:295 0.0349129
lASIG5V/1157 ASIG5V:2305 ASIG5V:263 402.919f 
rASIG5V/1158 ASIG5V:2305 ASIG5V:227 0.0349129
rASIG5V/1159 ASIG5V:227 X46/X28/D0:neg 0.445714
lASIG5V/1160 ASIG5V:2303 ASIG5V:225 136.992f 
rASIG5V/1161 ASIG5V:2303 ASIG5V:1308 0.0118704
lASIG5V/1162 ASIG5V:2301 ASIG5V:261 402.919f 
rASIG5V/1163 ASIG5V:2301 ASIG5V:225 0.0349129
rASIG5V/1164 ASIG5V:225 X46/X28/D0:neg 0.445714
lASIG5V/1165 ASIG5V:2299 ASIG5V:223 402.919f 
rASIG5V/1166 ASIG5V:2299 ASIG5V:291 0.0349129
lASIG5V/1167 ASIG5V:2297 ASIG5V:259 402.919f 
rASIG5V/1168 ASIG5V:2297 ASIG5V:223 0.0349129
rASIG5V/1169 ASIG5V:223 X46/X28/D0:neg 0.445714
lASIG5V/1170 ASIG5V:2295 ASIG5V:221 8.05837f 
rASIG5V/1171 ASIG5V:2295 ASIG5V:1292 0.000698258
lASIG5V/1172 ASIG5V:2293 ASIG5V:257 604.378f 
rASIG5V/1173 ASIG5V:2293 ASIG5V:221 0.0523694
rASIG5V/1174 ASIG5V:221 X46/X28/D0:neg 0.445714
lASIG5V/1175 ASIG5V:2291 ASIG5V:219 402.919f 
rASIG5V/1176 ASIG5V:2291 ASIG5V:287 0.0349129
lASIG5V/1177 ASIG5V:2289 ASIG5V:255 402.919f 
rASIG5V/1178 ASIG5V:2289 ASIG5V:219 0.0349129
rASIG5V/1179 ASIG5V:219 X46/X28/D0:neg 0.445714
lASIG5V/1180 ASIG5V:2287 ASIG5V:217 80.5837f 
rASIG5V/1181 ASIG5V:2287 ASIG5V:1276 0.00698258
lASIG5V/1182 ASIG5V:2285 ASIG5V:253 402.919f 
rASIG5V/1183 ASIG5V:2285 ASIG5V:217 0.0349129
rASIG5V/1184 ASIG5V:217 X46/X28/D0:neg 0.445714
lASIG5V/1185 ASIG5V:2283 ASIG5V:215 402.919f 
rASIG5V/1186 ASIG5V:2283 ASIG5V:283 0.0349129
lASIG5V/1187 ASIG5V:2281 ASIG5V:251 402.919f 
rASIG5V/1188 ASIG5V:2281 ASIG5V:215 0.0349129
rASIG5V/1189 ASIG5V:215 X46/X28/D0:neg 0.445714
lASIG5V/1190 ASIG5V:2279 ASIG5V:213 402.919f 
rASIG5V/1191 ASIG5V:2279 ASIG5V:281 0.0349129
lASIG5V/1192 ASIG5V:2277 ASIG5V:1260 48.3502f 
rASIG5V/1193 ASIG5V:2277 ASIG5V:213 0.00418955
rASIG5V/1194 ASIG5V:213 X46/X28/D0:neg 0.445714
rASIG5V/1195 X46/X27/D0:neg ASIG5V:1374 0.445714
lASIG5V/1196 ASIG5V:2275 ASIG5V:206 539.467f 
rASIG5V/1197 ASIG5V:2275 ASIG5V:1374 0.0470395
rASIG5V/1198 X46/X27/D0:neg ASIG5V:206 0.445714
rASIG5V/1199 X46/X27/D0:neg ASIG5V:204 0.445714
lASIG5V/1200 ASIG5V:2273 ASIG5V:202 370.047f 
rASIG5V/1201 ASIG5V:2273 ASIG5V:1358 0.0322668
rASIG5V/1202 X46/X27/D0:neg ASIG5V:202 0.445714
rASIG5V/1203 X46/X27/D0:neg ASIG5V:200 0.445714
lASIG5V/1204 ASIG5V:2271 ASIG5V:198 205.087f 
rASIG5V/1205 ASIG5V:2271 ASIG5V:1342 0.0178828
rASIG5V/1206 X46/X27/D0:neg ASIG5V:198 0.445714
rASIG5V/1207 X46/X27/D0:neg ASIG5V:196 0.445714
lASIG5V/1208 ASIG5V:2269 ASIG5V:194 285.338f 
rASIG5V/1209 ASIG5V:2269 ASIG5V:1326 0.0248804
rASIG5V/1210 X46/X27/D0:neg ASIG5V:194 0.445714
rASIG5V/1211 X46/X27/D0:neg ASIG5V:192 0.445714
rASIG5V/1212 ASIG5V:190 X46/X27/D0:neg 0.445714
lASIG5V/1213 ASIG5V:2267 ASIG5V:1310 294.255f 
rASIG5V/1214 ASIG5V:2267 ASIG5V:188 0.0256579
rASIG5V/1215 ASIG5V:188 X46/X27/D0:neg 0.445714
rASIG5V/1216 ASIG5V:186 X46/X27/D0:neg 0.445714
lASIG5V/1217 ASIG5V:2265 ASIG5V:1294 214.003f 
rASIG5V/1218 ASIG5V:2265 ASIG5V:184 0.0186603
rASIG5V/1219 ASIG5V:184 X46/X27/D0:neg 0.445714
rASIG5V/1220 ASIG5V:182 X46/X27/D0:neg 0.445714
lASIG5V/1221 ASIG5V:2263 ASIG5V:1278 356.672f 
rASIG5V/1222 ASIG5V:2263 ASIG5V:180 0.0311005
rASIG5V/1223 ASIG5V:180 X46/X27/D0:neg 0.445714
rASIG5V/1224 ASIG5V:178 X46/X27/D0:neg 0.445714
rASIG5V/1225 ASIG5V:176 X46/X27/D0:neg 0.445714
lASIG5V/1226 ASIG5V:2261 X46/X27/D0:neg 445.84f 
rASIG5V/1227 ASIG5V:2261 ASIG5V:176 0.23574
lASIG5V/1228 ASIG5V:2259 ASIG5V:204 450.299f 
rASIG5V/1229 ASIG5V:2259 ASIG5V:170 0.0392644
rASIG5V/1230 X46/X27/D0:neg ASIG5V:170 0.445714
lASIG5V/1231 ASIG5V:2257 ASIG5V:1358 80.2513f 
rASIG5V/1232 ASIG5V:2257 ASIG5V:168 0.00699761
rASIG5V/1233 X46/X27/D0:neg ASIG5V:168 0.445714
lASIG5V/1234 ASIG5V:2255 ASIG5V:200 450.299f 
rASIG5V/1235 ASIG5V:2255 ASIG5V:166 0.0392644
rASIG5V/1236 X46/X27/D0:neg ASIG5V:166 0.445714
lASIG5V/1237 ASIG5V:2253 ASIG5V:1342 17.8336f 
rASIG5V/1238 ASIG5V:2253 ASIG5V:164 0.00155502
rASIG5V/1239 X46/X27/D0:neg ASIG5V:164 0.445714
lASIG5V/1240 ASIG5V:2251 ASIG5V:196 445.84f 
rASIG5V/1241 ASIG5V:2251 ASIG5V:162 0.0388756
rASIG5V/1242 X46/X27/D0:neg ASIG5V:162 0.445714
lASIG5V/1243 ASIG5V:2249 ASIG5V:1326 160.503f 
rASIG5V/1244 ASIG5V:2249 ASIG5V:160 0.0139952
rASIG5V/1245 X46/X27/D0:neg ASIG5V:160 0.445714
lASIG5V/1246 ASIG5V:2247 ASIG5V:192 445.84f 
rASIG5V/1247 ASIG5V:2247 ASIG5V:158 0.0388756
rASIG5V/1248 X46/X27/D0:neg ASIG5V:158 0.445714
lASIG5V/1249 ASIG5V:2245 ASIG5V:190 445.84f 
rASIG5V/1250 ASIG5V:2245 ASIG5V:156 0.0388756
rASIG5V/1251 ASIG5V:156 X46/X27/D0:neg 0.445714
lASIG5V/1252 ASIG5V:2243 ASIG5V:188 445.84f 
rASIG5V/1253 ASIG5V:2243 ASIG5V:154 0.0388756
rASIG5V/1254 ASIG5V:154 X46/X27/D0:neg 0.445714
lASIG5V/1255 ASIG5V:2241 ASIG5V:186 222.92f 
rASIG5V/1256 ASIG5V:2241 ASIG5V:152 0.0194378
rASIG5V/1257 ASIG5V:152 X46/X27/D0:neg 0.445714
lASIG5V/1258 ASIG5V:2239 ASIG5V:184 445.84f 
rASIG5V/1259 ASIG5V:2239 ASIG5V:150 0.0388756
rASIG5V/1260 ASIG5V:150 X46/X27/D0:neg 0.445714
lASIG5V/1261 ASIG5V:2237 ASIG5V:182 445.84f 
rASIG5V/1262 ASIG5V:2237 ASIG5V:148 0.0388756
rASIG5V/1263 ASIG5V:148 X46/X27/D0:neg 0.445714
lASIG5V/1264 ASIG5V:2235 ASIG5V:180 445.84f 
rASIG5V/1265 ASIG5V:2235 ASIG5V:146 0.0388756
rASIG5V/1266 ASIG5V:146 X46/X27/D0:neg 0.445714
lASIG5V/1267 ASIG5V:2233 ASIG5V:144 392.339f 
rASIG5V/1268 ASIG5V:2233 ASIG5V:1262 0.0342105
lASIG5V/1269 ASIG5V:2231 ASIG5V:178 445.84f 
rASIG5V/1270 ASIG5V:2231 ASIG5V:144 0.0388756
rASIG5V/1271 ASIG5V:144 X46/X27/D0:neg 0.445714
lASIG5V/1272 ASIG5V:2229 ASIG5V:138 450.299f 
rASIG5V/1273 ASIG5V:2229 ASIG5V:206 0.0392644
lASIG5V/1274 ASIG5V:2227 ASIG5V:138 450.299f 
rASIG5V/1275 ASIG5V:2227 X46/X27/D0:neg 0.271523
rASIG5V/1276 X46/X27/D0:neg ASIG5V:138 0.445714
lASIG5V/1277 ASIG5V:2225 ASIG5V:136 450.299f 
rASIG5V/1278 ASIG5V:2225 ASIG5V:204 0.0392644
lASIG5V/1279 ASIG5V:2223 ASIG5V:1374 361.131f 
rASIG5V/1280 ASIG5V:2223 ASIG5V:136 0.0314892
rASIG5V/1281 X46/X27/D0:neg ASIG5V:136 0.445714
lASIG5V/1282 ASIG5V:2221 ASIG5V:134 450.299f 
rASIG5V/1283 ASIG5V:2221 ASIG5V:202 0.0392644
lASIG5V/1284 ASIG5V:2219 ASIG5V:170 450.299f 
rASIG5V/1285 ASIG5V:2219 ASIG5V:134 0.0392644
rASIG5V/1286 X46/X27/D0:neg ASIG5V:134 0.445714
lASIG5V/1287 ASIG5V:2217 ASIG5V:132 450.299f 
rASIG5V/1288 ASIG5V:2217 ASIG5V:200 0.0392644
lASIG5V/1289 ASIG5V:2215 ASIG5V:168 450.299f 
rASIG5V/1290 ASIG5V:2215 ASIG5V:132 0.0392644
rASIG5V/1291 X46/X27/D0:neg ASIG5V:132 0.445714
lASIG5V/1292 ASIG5V:2213 ASIG5V:130 445.84f 
rASIG5V/1293 ASIG5V:2213 ASIG5V:198 0.0388756
lASIG5V/1294 ASIG5V:2211 ASIG5V:166 450.299f 
rASIG5V/1295 ASIG5V:2211 ASIG5V:130 0.0392644
rASIG5V/1296 X46/X27/D0:neg ASIG5V:130 0.445714
lASIG5V/1297 ASIG5V:2209 ASIG5V:128 222.92f 
rASIG5V/1298 ASIG5V:2209 ASIG5V:196 0.0194378
lASIG5V/1299 ASIG5V:2207 ASIG5V:164 668.761f 
rASIG5V/1300 ASIG5V:2207 ASIG5V:128 0.0583134
rASIG5V/1301 X46/X27/D0:neg ASIG5V:128 0.445714
lASIG5V/1302 ASIG5V:2205 ASIG5V:126 445.84f 
rASIG5V/1303 ASIG5V:2205 ASIG5V:194 0.0388756
lASIG5V/1304 ASIG5V:2203 ASIG5V:162 445.84f 
rASIG5V/1305 ASIG5V:2203 ASIG5V:126 0.0388756
rASIG5V/1306 X46/X27/D0:neg ASIG5V:126 0.445714
lASIG5V/1307 ASIG5V:2201 ASIG5V:124 445.84f 
rASIG5V/1308 ASIG5V:2201 ASIG5V:192 0.0388756
lASIG5V/1309 ASIG5V:2199 ASIG5V:160 445.84f 
rASIG5V/1310 ASIG5V:2199 ASIG5V:124 0.0388756
rASIG5V/1311 X46/X27/D0:neg ASIG5V:124 0.445714
lASIG5V/1312 ASIG5V:2197 ASIG5V:122 445.84f 
rASIG5V/1313 ASIG5V:2197 ASIG5V:190 0.0388756
lASIG5V/1314 ASIG5V:2195 ASIG5V:158 445.84f 
rASIG5V/1315 ASIG5V:2195 ASIG5V:122 0.0388756
rASIG5V/1316 ASIG5V:122 X46/X27/D0:neg 0.445714
lASIG5V/1317 ASIG5V:2193 ASIG5V:120 151.586f 
rASIG5V/1318 ASIG5V:2193 ASIG5V:1310 0.0132177
lASIG5V/1319 ASIG5V:2191 ASIG5V:156 445.84f 
rASIG5V/1320 ASIG5V:2191 ASIG5V:120 0.0388756
rASIG5V/1321 ASIG5V:120 X46/X27/D0:neg 0.445714
lASIG5V/1322 ASIG5V:2189 ASIG5V:118 445.84f 
rASIG5V/1323 ASIG5V:2189 ASIG5V:186 0.0388756
lASIG5V/1324 ASIG5V:2187 ASIG5V:154 445.84f 
rASIG5V/1325 ASIG5V:2187 ASIG5V:118 0.0388756
rASIG5V/1326 ASIG5V:118 X46/X27/D0:neg 0.445714
lASIG5V/1327 ASIG5V:2185 ASIG5V:116 8.91681f 
rASIG5V/1328 ASIG5V:2185 ASIG5V:1294 0.000777512
lASIG5V/1329 ASIG5V:2183 ASIG5V:152 668.761f 
rASIG5V/1330 ASIG5V:2183 ASIG5V:116 0.0583134
rASIG5V/1331 ASIG5V:116 X46/X27/D0:neg 0.445714
lASIG5V/1332 ASIG5V:2181 ASIG5V:114 445.84f 
rASIG5V/1333 ASIG5V:2181 ASIG5V:182 0.0388756
lASIG5V/1334 ASIG5V:2179 ASIG5V:150 445.84f 
rASIG5V/1335 ASIG5V:2179 ASIG5V:114 0.0388756
rASIG5V/1336 ASIG5V:114 X46/X27/D0:neg 0.445714
lASIG5V/1337 ASIG5V:2177 ASIG5V:112 89.1681f 
rASIG5V/1338 ASIG5V:2177 ASIG5V:1278 0.00777512
lASIG5V/1339 ASIG5V:2175 ASIG5V:148 445.84f 
rASIG5V/1340 ASIG5V:2175 ASIG5V:112 0.0388756
rASIG5V/1341 ASIG5V:112 X46/X27/D0:neg 0.445714
lASIG5V/1342 ASIG5V:2173 ASIG5V:110 445.84f 
rASIG5V/1343 ASIG5V:2173 ASIG5V:178 0.0388756
lASIG5V/1344 ASIG5V:2171 ASIG5V:146 445.84f 
rASIG5V/1345 ASIG5V:2171 ASIG5V:110 0.0388756
rASIG5V/1346 ASIG5V:110 X46/X27/D0:neg 0.445714
lASIG5V/1347 ASIG5V:2169 ASIG5V:108 445.84f 
rASIG5V/1348 ASIG5V:2169 ASIG5V:176 0.0388756
lASIG5V/1349 ASIG5V:2167 ASIG5V:1262 53.5008f 
rASIG5V/1350 ASIG5V:2167 ASIG5V:108 0.00466507
rASIG5V/1351 ASIG5V:108 X46/X27/D0:neg 0.445714
rASIG5V/1352 X46/X26/D0:neg ASIG5V:1376 0.445714
lASIG5V/1353 ASIG5V:2165 ASIG5V:101 565.99f 
rASIG5V/1354 ASIG5V:2165 ASIG5V:1376 0.0498351
rASIG5V/1355 X46/X26/D0:neg ASIG5V:101 0.445714
rASIG5V/1356 X46/X26/D0:neg ASIG5V:99 0.445714
lASIG5V/1357 ASIG5V:2163 ASIG5V:97 388.241f 
rASIG5V/1358 ASIG5V:2163 ASIG5V:1360 0.0341844
rASIG5V/1359 X46/X26/D0:neg ASIG5V:97 0.445714
rASIG5V/1360 X46/X26/D0:neg ASIG5V:95 0.445714
lASIG5V/1361 ASIG5V:2161 ASIG5V:93 215.17f 
rASIG5V/1362 ASIG5V:2161 ASIG5V:1344 0.0189456
rASIG5V/1363 X46/X26/D0:neg ASIG5V:93 0.445714
rASIG5V/1364 X46/X26/D0:neg ASIG5V:91 0.445714
lASIG5V/1365 ASIG5V:2159 ASIG5V:89 299.367f 
rASIG5V/1366 ASIG5V:2159 ASIG5V:1328 0.026359
rASIG5V/1367 X46/X26/D0:neg ASIG5V:89 0.445714
rASIG5V/1368 X46/X26/D0:neg ASIG5V:87 0.445714
rASIG5V/1369 ASIG5V:85 X46/X26/D0:neg 0.445714
lASIG5V/1370 ASIG5V:2157 ASIG5V:1312 308.722f 
rASIG5V/1371 ASIG5V:2157 ASIG5V:83 0.0271828
rASIG5V/1372 ASIG5V:83 X46/X26/D0:neg 0.445714
rASIG5V/1373 ASIG5V:81 X46/X26/D0:neg 0.445714
lASIG5V/1374 ASIG5V:2155 ASIG5V:1296 224.525f 
rASIG5V/1375 ASIG5V:2155 ASIG5V:79 0.0197693
rASIG5V/1376 ASIG5V:79 X46/X26/D0:neg 0.445714
rASIG5V/1377 ASIG5V:77 X46/X26/D0:neg 0.445714
lASIG5V/1378 ASIG5V:2153 ASIG5V:1280 374.209f 
rASIG5V/1379 ASIG5V:2153 ASIG5V:75 0.0329488
rASIG5V/1380 ASIG5V:75 X46/X26/D0:neg 0.445714
rASIG5V/1381 ASIG5V:73 X46/X26/D0:neg 0.445714
rASIG5V/1382 ASIG5V:71 X46/X26/D0:neg 0.445714
lASIG5V/1383 ASIG5V:2151 X46/X26/D0:neg 467.761f 
rASIG5V/1384 ASIG5V:2151 ASIG5V:71 0.2388
lASIG5V/1385 ASIG5V:2149 ASIG5V:99 472.438f 
rASIG5V/1386 ASIG5V:2149 ASIG5V:65 0.0415979
rASIG5V/1387 X46/X26/D0:neg ASIG5V:65 0.445714
lASIG5V/1388 ASIG5V:2147 ASIG5V:1360 84.1969f 
rASIG5V/1389 ASIG5V:2147 ASIG5V:63 0.00741348
rASIG5V/1390 X46/X26/D0:neg ASIG5V:63 0.445714
lASIG5V/1391 ASIG5V:2145 ASIG5V:95 472.438f 
rASIG5V/1392 ASIG5V:2145 ASIG5V:61 0.0415979
rASIG5V/1393 X46/X26/D0:neg ASIG5V:61 0.445714
lASIG5V/1394 ASIG5V:2143 ASIG5V:1344 18.7104f 
rASIG5V/1395 ASIG5V:2143 ASIG5V:59 0.00164744
rASIG5V/1396 X46/X26/D0:neg ASIG5V:59 0.445714
lASIG5V/1397 ASIG5V:2141 ASIG5V:91 467.761f 
rASIG5V/1398 ASIG5V:2141 ASIG5V:57 0.041186
rASIG5V/1399 X46/X26/D0:neg ASIG5V:57 0.445714
lASIG5V/1400 ASIG5V:2139 ASIG5V:1328 168.394f 
rASIG5V/1401 ASIG5V:2139 ASIG5V:55 0.014827
rASIG5V/1402 X46/X26/D0:neg ASIG5V:55 0.445714
lASIG5V/1403 ASIG5V:2137 ASIG5V:87 467.761f 
rASIG5V/1404 ASIG5V:2137 ASIG5V:53 0.041186
rASIG5V/1405 X46/X26/D0:neg ASIG5V:53 0.445714
lASIG5V/1406 ASIG5V:2135 ASIG5V:85 467.761f 
rASIG5V/1407 ASIG5V:2135 ASIG5V:51 0.041186
rASIG5V/1408 ASIG5V:51 X46/X26/D0:neg 0.445714
lASIG5V/1409 ASIG5V:2133 ASIG5V:83 467.761f 
rASIG5V/1410 ASIG5V:2133 ASIG5V:49 0.041186
rASIG5V/1411 ASIG5V:49 X46/X26/D0:neg 0.445714
lASIG5V/1412 ASIG5V:2131 ASIG5V:81 233.88f 
rASIG5V/1413 ASIG5V:2131 ASIG5V:47 0.020593
rASIG5V/1414 ASIG5V:47 X46/X26/D0:neg 0.445714
lASIG5V/1415 ASIG5V:2129 ASIG5V:79 467.761f 
rASIG5V/1416 ASIG5V:2129 ASIG5V:45 0.041186
rASIG5V/1417 ASIG5V:45 X46/X26/D0:neg 0.445714
lASIG5V/1418 ASIG5V:2127 ASIG5V:77 467.761f 
rASIG5V/1419 ASIG5V:2127 ASIG5V:43 0.041186
rASIG5V/1420 ASIG5V:43 X46/X26/D0:neg 0.445714
lASIG5V/1421 ASIG5V:2125 ASIG5V:75 467.761f 
rASIG5V/1422 ASIG5V:2125 ASIG5V:41 0.041186
rASIG5V/1423 ASIG5V:41 X46/X26/D0:neg 0.445714
lASIG5V/1424 ASIG5V:2123 ASIG5V:39 411.629f 
rASIG5V/1425 ASIG5V:2123 ASIG5V:1264 0.0362437
lASIG5V/1426 ASIG5V:2121 ASIG5V:73 467.761f 
rASIG5V/1427 ASIG5V:2121 ASIG5V:39 0.041186
rASIG5V/1428 ASIG5V:39 X46/X26/D0:neg 0.445714
lASIG5V/1429 ASIG5V:2119 ASIG5V:33 472.438f 
rASIG5V/1430 ASIG5V:2119 ASIG5V:101 0.0415979
lASIG5V/1431 ASIG5V:2117 ASIG5V:33 472.438f 
rASIG5V/1432 ASIG5V:2117 X46/X26/D0:neg 0.274391
rASIG5V/1433 X46/X26/D0:neg ASIG5V:33 0.445714
lASIG5V/1434 ASIG5V:2115 ASIG5V:31 472.438f 
rASIG5V/1435 ASIG5V:2115 ASIG5V:99 0.0415979
lASIG5V/1436 ASIG5V:2113 ASIG5V:1376 378.886f 
rASIG5V/1437 ASIG5V:2113 ASIG5V:31 0.0333607
rASIG5V/1438 X46/X26/D0:neg ASIG5V:31 0.445714
lASIG5V/1439 ASIG5V:2111 ASIG5V:29 472.438f 
rASIG5V/1440 ASIG5V:2111 ASIG5V:97 0.0415979
lASIG5V/1441 ASIG5V:2109 ASIG5V:65 472.438f 
rASIG5V/1442 ASIG5V:2109 ASIG5V:29 0.0415979
rASIG5V/1443 X46/X26/D0:neg ASIG5V:29 0.445714
lASIG5V/1444 ASIG5V:2107 ASIG5V:27 472.438f 
rASIG5V/1445 ASIG5V:2107 ASIG5V:95 0.0415979
lASIG5V/1446 ASIG5V:2105 ASIG5V:63 472.438f 
rASIG5V/1447 ASIG5V:2105 ASIG5V:27 0.0415979
rASIG5V/1448 X46/X26/D0:neg ASIG5V:27 0.445714
lASIG5V/1449 ASIG5V:2103 ASIG5V:25 467.761f 
rASIG5V/1450 ASIG5V:2103 ASIG5V:93 0.041186
lASIG5V/1451 ASIG5V:2101 ASIG5V:61 472.438f 
rASIG5V/1452 ASIG5V:2101 ASIG5V:25 0.0415979
rASIG5V/1453 X46/X26/D0:neg ASIG5V:25 0.445714
lASIG5V/1454 ASIG5V:2099 ASIG5V:23 233.88f 
rASIG5V/1455 ASIG5V:2099 ASIG5V:91 0.020593
lASIG5V/1456 ASIG5V:2097 ASIG5V:59 701.641f 
rASIG5V/1457 ASIG5V:2097 ASIG5V:23 0.061779
rASIG5V/1458 X46/X26/D0:neg ASIG5V:23 0.445714
lASIG5V/1459 ASIG5V:2095 ASIG5V:21 467.761f 
rASIG5V/1460 ASIG5V:2095 ASIG5V:89 0.041186
lASIG5V/1461 ASIG5V:2093 ASIG5V:57 467.761f 
rASIG5V/1462 ASIG5V:2093 ASIG5V:21 0.041186
rASIG5V/1463 X46/X26/D0:neg ASIG5V:21 0.445714
lASIG5V/1464 ASIG5V:2091 ASIG5V:19 467.761f 
rASIG5V/1465 ASIG5V:2091 ASIG5V:87 0.041186
lASIG5V/1466 ASIG5V:2089 ASIG5V:55 467.761f 
rASIG5V/1467 ASIG5V:2089 ASIG5V:19 0.041186
rASIG5V/1468 X46/X26/D0:neg ASIG5V:19 0.445714
lASIG5V/1469 ASIG5V:2087 ASIG5V:17 467.761f 
rASIG5V/1470 ASIG5V:2087 ASIG5V:85 0.041186
lASIG5V/1471 ASIG5V:2085 ASIG5V:53 467.761f 
rASIG5V/1472 ASIG5V:2085 ASIG5V:17 0.041186
rASIG5V/1473 ASIG5V:17 X46/X26/D0:neg 0.445714
lASIG5V/1474 ASIG5V:2083 ASIG5V:15 159.039f 
rASIG5V/1475 ASIG5V:2083 ASIG5V:1312 0.0140032
lASIG5V/1476 ASIG5V:2081 ASIG5V:51 467.761f 
rASIG5V/1477 ASIG5V:2081 ASIG5V:15 0.041186
rASIG5V/1478 ASIG5V:15 X46/X26/D0:neg 0.445714
lASIG5V/1479 ASIG5V:2079 ASIG5V:13 467.761f 
rASIG5V/1480 ASIG5V:2079 ASIG5V:81 0.041186
lASIG5V/1481 ASIG5V:2077 ASIG5V:49 467.761f 
rASIG5V/1482 ASIG5V:2077 ASIG5V:13 0.041186
rASIG5V/1483 ASIG5V:13 X46/X26/D0:neg 0.445714
lASIG5V/1484 ASIG5V:2075 ASIG5V:11 9.35521f 
rASIG5V/1485 ASIG5V:2075 ASIG5V:1296 0.00082372
lASIG5V/1486 ASIG5V:2073 ASIG5V:47 701.641f 
rASIG5V/1487 ASIG5V:2073 ASIG5V:11 0.061779
rASIG5V/1488 ASIG5V:11 X46/X26/D0:neg 0.445714
lASIG5V/1489 ASIG5V:2071 ASIG5V:9 467.761f 
rASIG5V/1490 ASIG5V:2071 ASIG5V:77 0.041186
lASIG5V/1491 ASIG5V:2069 ASIG5V:45 467.761f 
rASIG5V/1492 ASIG5V:2069 ASIG5V:9 0.041186
rASIG5V/1493 ASIG5V:9 X46/X26/D0:neg 0.445714
lASIG5V/1494 ASIG5V:2067 ASIG5V:7 93.5521f 
rASIG5V/1495 ASIG5V:2067 ASIG5V:1280 0.0082372
lASIG5V/1496 ASIG5V:2065 ASIG5V:43 467.761f 
rASIG5V/1497 ASIG5V:2065 ASIG5V:7 0.041186
rASIG5V/1498 ASIG5V:7 X46/X26/D0:neg 0.445714
lASIG5V/1499 ASIG5V:2063 ASIG5V:5 467.761f 
rASIG5V/1500 ASIG5V:2063 ASIG5V:73 0.041186
lASIG5V/1501 ASIG5V:2061 ASIG5V:41 467.761f 
rASIG5V/1502 ASIG5V:2061 ASIG5V:5 0.041186
rASIG5V/1503 ASIG5V:5 X46/X26/D0:neg 0.445714
lASIG5V/1504 ASIG5V:2059 ASIG5V:3 467.761f 
rASIG5V/1505 ASIG5V:2059 ASIG5V:71 0.041186
lASIG5V/1506 ASIG5V:2057 ASIG5V:1264 56.1313f 
rASIG5V/1507 ASIG5V:2057 ASIG5V:3 0.00494232
rASIG5V/1508 ASIG5V:3 X46/X26/D0:neg 0.445714
XR0 R0:pos R0:neg rm2 r_width=2.54e-06 r_length=2.76e-07
XR1 R1:pos R1:neg rm2 r_width=2.54e-06 r_length=2.76e-07
XR2 R2:pos R2:neg rm2 r_width=2.54e-06 r_length=2.76e-07
XR3 R3:pos R3:neg rm2 r_width=2.54e-06 r_length=2.76e-07
XR4 R4:pos R4:neg rm2 r_width=2.54e-06 r_length=2.76e-07
XR5 R5:pos R5:neg rm2 r_width=2.54e-06 r_length=2.76e-07
XR6 R6:pos R6:neg rm2 r_width=2.54e-06 r_length=2.76e-07
XR7 R7:pos R7:neg rm2 r_width=2.54e-06 r_length=2.76e-07
dX27/D0 DVSS X27/D0:neg diode_nd2ps_06v0  area=4e-11 pj=8.2e-05 M=1
dX28/D0 DVSS X28/D0:neg diode_nd2ps_06v0  area=4e-11 pj=8.2e-05 M=1
dX29/D0 DVSS X29/D0:neg diode_nd2ps_06v0  area=4e-11 pj=8.2e-05 M=1
dX30/D0 DVSS X30/D0:neg diode_nd2ps_06v0  area=4e-11 pj=8.2e-05 M=1
dX46/X26/D0 DVSS X46/X26/D0:neg diode_nd2ps_06v0  area=1.5e-10 pj=0.000106 M=1
dX46/X27/D0 DVSS X46/X27/D0:neg diode_nd2ps_06v0  area=1.5e-10 pj=0.000106 M=1
dX46/X28/D0 DVSS X46/X28/D0:neg diode_nd2ps_06v0  area=1.5e-10 pj=0.000106 M=1
dX46/X29/D0 DVSS X46/X29/D0:neg diode_nd2ps_06v0  area=1.5e-10 pj=0.000106 M=1
dX46/X30/D0 X46/X30/D0:pos X46/X30/D0:neg diode_pd2nw_06v0  area=1.5e-10 pj=0.000106 M=1
dX46/X31/D0 X46/X31/D0:pos X46/X31/D0:neg diode_pd2nw_06v0  area=1.5e-10 pj=0.000106 M=1
dX46/X32/D0 X46/X32/D0:pos X46/X32/D0:neg diode_pd2nw_06v0  area=1.5e-10 pj=0.000106 M=1
dX46/X33/D0 X46/X33/D0:pos X46/X33/D0:neg diode_pd2nw_06v0  area=1.5e-10 pj=0.000106 M=1
XX48/X1/X0/C0 X48/X1/X0/C0:pos DVSS cap_nmos_06v0        c_length=1.5e-05 c_width=1.5e-05
XX48/X1/X1/C0 X48/X1/X1/C0:pos DVSS cap_nmos_06v0        c_length=1.5e-05 c_width=1.5e-05
XX48/X2/X0/C0 X48/X2/X0/C0:pos DVSS cap_nmos_06v0        c_length=1.5e-05 c_width=1.5e-05
XX48/X2/X1/C0 X48/X2/X1/C0:pos DVSS cap_nmos_06v0        c_length=1.5e-05 c_width=1.5e-05
XX49/X0/X1/X0/C0 X49/X0/X1/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX49/X0/X1/X1/C0 X49/X0/X1/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX49/X0/X2/X0/C0 X49/X0/X2/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX49/X0/X2/X1/C0 X49/X0/X2/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX49/X1/X1/X0/C0 X49/X1/X1/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX49/X1/X1/X1/C0 X49/X1/X1/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX49/X1/X2/X0/C0 X49/X1/X2/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX49/X1/X2/X1/C0 X49/X1/X2/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX50/X0/X1/X0/C0 X50/X0/X1/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX50/X0/X1/X1/C0 X50/X0/X1/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX50/X0/X2/X0/C0 X50/X0/X2/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX50/X0/X2/X1/C0 X50/X0/X2/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX50/X1/X1/X0/C0 X50/X1/X1/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX50/X1/X1/X1/C0 X50/X1/X1/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX50/X1/X2/X0/C0 X50/X1/X2/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX50/X1/X2/X1/C0 X50/X1/X2/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX51/X0/X1/X0/C0 X51/X0/X1/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX51/X0/X1/X1/C0 X51/X0/X1/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX51/X0/X2/X0/C0 X51/X0/X2/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX51/X0/X2/X1/C0 X51/X0/X2/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX51/X1/X1/X0/C0 X51/X1/X1/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX51/X1/X1/X1/C0 X51/X1/X1/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX51/X1/X2/X0/C0 X51/X1/X2/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX51/X1/X2/X1/C0 X51/X1/X2/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX52/X0/X1/X0/C0 X52/X0/X1/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX52/X0/X1/X1/C0 X52/X0/X1/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX52/X0/X2/X0/C0 X52/X0/X2/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX52/X0/X2/X1/C0 X52/X0/X2/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX52/X1/X1/X0/C0 X52/X1/X1/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX52/X1/X1/X1/C0 X52/X1/X1/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX52/X1/X2/X0/C0 X52/X1/X2/X0/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
XX52/X1/X2/X1/C0 X52/X1/X2/X1/C0:pos DVSS cap_nmos_06v0  c_length=1.5e-05 c_width=1.5e-05
.ends
